# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0050 ;

LAYER poly
  TYPE CUT ;
  SPACING 0.072 ;
END poly

LAYER active
  TYPE CUT ;
  SPACING 0.072 ;
END active

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.14 ;
  AREA 0.020000 ;
  WIDTH 0.070 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0    0.06 
	WIDTH 0.1  0.1 
	WIDTH 0.75 0.25 
	WIDTH 1.5  0.45 ; 
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.080 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.19 ;
  AREA 0.020000 ;
  WIDTH 0.070 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0.00 0.07 
	WIDTH 0.09 0.07 
	WIDTH 0.27 0.07 
	WIDTH 0.50 0.07 
	WIDTH 0.90 0.07 
	WIDTH 1.50 0.07 ;
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.090 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.14 ;
  AREA 0.020000 ;
  WIDTH 0.070 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0.00 0.07 
	WIDTH 0.09 0.07 
	WIDTH 0.27 0.07 
	WIDTH 0.50 0.07 
	WIDTH 0.90 0.07 
	WIDTH 1.50 0.07 ;
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.090 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.28 ;
  AREA 0.020000 ;
  WIDTH 0.140 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0.00 0.14 
	WIDTH 0.27 0.14 
	WIDTH 0.50 0.14 
	WIDTH 0.90 0.14 
	WIDTH 1.50 0.14 ;
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.160 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.28 ;
  AREA 0.020000 ;
  WIDTH 0.140 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0.00 0.14 
	WIDTH 0.27 0.14 
	WIDTH 0.50 0.14 
	WIDTH 0.90 0.14 
	WIDTH 1.50 0.14 ;
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal5

LAYER via5
  TYPE CUT ;
  SPACING 0.160 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.28 ;
  AREA 0.020000 ;
  WIDTH 0.140 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0.00 0.14 
	WIDTH 0.27 0.14 
	WIDTH 0.50 0.14 
	WIDTH 0.90 0.14 
	WIDTH 1.50 0.14 ;
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal6

LAYER via6
  TYPE CUT ;
  SPACING 0.160 ;
END via6

LAYER metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.80 ;
  AREA 0.020000 ;
  WIDTH 0.400 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0.00 0.40 
	WIDTH 0.50 0.40 
	WIDTH 0.90 0.40 
	WIDTH 1.50 0.40 ;
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal7

LAYER via7
  TYPE CUT ;
  SPACING 0.440 ;
END via7

LAYER metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.80 ;
  AREA 0.020000 ;
  WIDTH 0.400 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0.00 0.40 
	WIDTH 0.50 0.40 
	WIDTH 0.90 0.40 
	WIDTH 1.50 0.40 ;
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal8

LAYER via8
  TYPE CUT ;
  SPACING 0.440 ;
END via8

LAYER metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.60 ;
  AREA 0.020000 ;
  WIDTH 0.800 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0.00 0.80 
	WIDTH 0.90 0.80 
	WIDTH 1.50 0.80 ;
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal9

LAYER via9
  TYPE CUT ;
  SPACING 0.880 ;
END via9

LAYER metal10
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.60 ;
  AREA 0.020000 ;
  WIDTH 0.800 ;
  SPACINGTABLE
	PARALLELRUNLENGTH 0
	WIDTH 0.00 0.80 
	WIDTH 0.90 0.80 
	WIDTH 1.50 0.80 ;
  SPACING 0.09 ENDOFLINE 0.09 WITHIN 0.025 ;
END metal10

LAYER OVERLAP
  TYPE CUT ;
  SPACING 0.072 ;
END OVERLAP

