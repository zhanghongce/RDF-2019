module ac97_ctrl (
	x977,
	x96,
	x940,
	x906,
	x889,
	x868,
	x84,
	x837,
	x821,
	x806,
	x786,
	x77,
	x765,
	x744,
	x718,
	x699,
	x681,
	x657,
	x638,
	x63,
	x620,
	x589,
	x561,
	x538,
	x522,
	x494,
	x476,
	x447,
	x420,
	x397,
	x390,
	x38,
	x379,
	x361,
	x342,
	x315,
	x30,
	x287,
	x264,
	x249,
	x234,
	x217,
	x195,
	x187,
	x1822,
	x179,
	x172,
	x1595,
	x1587,
	x1580,
	x1572,
	x1564,
	x1557,
	x1550,
	x1542,
	x1534,
	x1527,
	x1519,
	x1511,
	x1501,
	x1494,
	x149,
	x1486,
	x1479,
	x1467,
	x1459,
	x1451,
	x145,
	x1443,
	x1432,
	x1424,
	x1417,
	x1406,
	x14,
	x1398,
	x1390,
	x1382,
	x138,
	x1374,
	x1366,
	x1358,
	x1351,
	x1345,
	x1322,
	x131,
	x130657,
	x130656,
	x130655,
	x130654,
	x130653,
	x130652,
	x130651,
	x130650,
	x130649,
	x130648,
	x130647,
	x130646,
	x130645,
	x130644,
	x130643,
	x130642,
	x130641,
	x130640,
	x130639,
	x130638,
	x130637,
	x130636,
	x130635,
	x130634,
	x130633,
	x130632,
	x130631,
	x130630,
	x130629,
	x1286,
	x1261,
	x124,
	x1231,
	x1215,
	x1209,
	x1203,
	x1193,
	x1155,
	x114,
	x1126,
	x1101,
	x1062,
	x106,
	x1034,
	x101,
	x1006,
	x0,
	clk);
   input x977;
   output x96;
   input x940;
   input x906;
   input x889;
   input x868;
   output x84;
   input x837;
   input x821;
   input x806;
   output x786;
   output x77;
   output x765;
   output x744;
   output x718;
   output x699;
   output x681;
   output x657;
   output x638;
   output x63;
   output x620;
   output x589;
   output x561;
   output x538;
   output x522;
   output x494;
   output x476;
   output x447;
   output x420;
   output x397;
   output x390;
   output x38;
   output x379;
   output x361;
   output x342;
   output x315;
   output x30;
   output x287;
   output x264;
   output x249;
   output x234;
   output x217;
   output x195;
   output x187;
   input x1822;
   output x179;
   output x172;
   input x1595;
   input x1587;
   input x1580;
   input x1572;
   input x1564;
   input x1557;
   input x1550;
   input x1542;
   input x1534;
   input x1527;
   input x1519;
   input x1511;
   input x1501;
   input x1494;
   output x149;
   input x1486;
   input x1479;
   input x1467;
   input x1459;
   input x1451;
   output x145;
   input x1443;
   input x1432;
   input x1424;
   input x1417;
   input x1406;
   output x14;
   input x1398;
   input x1390;
   input x1382;
   output x138;
   input x1374;
   input x1366;
   input x1358;
   input x1351;
   input x1345;
   input x1322;
   output x131;
   input x130657;
   input x130656;
   input x130655;
   input x130654;
   input x130653;
   input x130652;
   input x130651;
   input x130650;
   input x130649;
   input x130648;
   input x130647;
   input x130646;
   input x130645;
   input x130644;
   input x130643;
   input x130642;
   input x130641;
   input x130640;
   input x130639;
   input x130638;
   input x130637;
   input x130636;
   input x130635;
   input x130634;
   input x130633;
   input x130632;
   input x130631;
   input x130630;
   input x130629;
   input x1286;
   input x1261;
   output x124;
   input x1231;
   input x1215;
   input x1209;
   input x1203;
   input x1193;
   input x1155;
   output x114;
   input x1126;
   input x1101;
   input x1062;
   output x106;
   input x1034;
   output x101;
   input x1006;
   output x0;
   input clk;

   // Internal wires
   wire x977;
   wire x96;
   wire x940;
   wire x906;
   wire x889;
   wire x868;
   wire x84;
   wire x837;
   wire x821;
   wire x806;
   wire x786;
   wire x77;
   wire x765;
   wire x744;
   wire x718;
   wire x699;
   wire x681;
   wire x657;
   wire x638;
   wire x63;
   wire x620;
   wire x589;
   wire x561;
   wire x538;
   wire x522;
   wire x494;
   wire x476;
   wire x447;
   wire x420;
   wire x397;
   wire x390;
   wire x38;
   wire x379;
   wire x361;
   wire x342;
   wire x315;
   wire x30;
   wire x287;
   wire x264;
   wire x249;
   wire x234;
   wire x217;
   wire x195;
   wire x187;
   wire x1822;
   wire x179;
   wire x172;
   wire x1595;
   wire x1587;
   wire x1580;
   wire x1572;
   wire x1564;
   wire x1557;
   wire x1550;
   wire x1542;
   wire x1534;
   wire x1527;
   wire x1519;
   wire x1511;
   wire x1501;
   wire x1494;
   wire x149;
   wire x1486;
   wire x1479;
   wire x1467;
   wire x1459;
   wire x1451;
   wire x145;
   wire x1443;
   wire x1432;
   wire x1424;
   wire x1417;
   wire x1406;
   wire x14;
   wire x1398;
   wire x1390;
   wire x1382;
   wire x138;
   wire x1374;
   wire x1366;
   wire x1358;
   wire x1351;
   wire x1345;
   wire x1322;
   wire x131;
   wire x130657;
   wire x130656;
   wire x130655;
   wire x130654;
   wire x130653;
   wire x130652;
   wire x130651;
   wire x130650;
   wire x130649;
   wire x130648;
   wire x130647;
   wire x130646;
   wire x130645;
   wire x130644;
   wire x130643;
   wire x130642;
   wire x130641;
   wire x130640;
   wire x130639;
   wire x130638;
   wire x130637;
   wire x130636;
   wire x130635;
   wire x130634;
   wire x130633;
   wire x130632;
   wire x130631;
   wire x130630;
   wire x130629;
   wire x1286;
   wire x1261;
   wire x124;
   wire x1231;
   wire x1215;
   wire x1209;
   wire x1203;
   wire x1193;
   wire x1155;
   wire x114;
   wire x1126;
   wire x1101;
   wire x1062;
   wire x106;
   wire x1034;
   wire x101;
   wire x1006;
   wire x0;
   wire new_n9999_;
   wire new_n9998_;
   wire new_n9997_1_;
   wire new_n9996_;
   wire new_n9995_;
   wire new_n9994_;
   wire new_n9993_;
   wire new_n9992_1_;
   wire new_n9991_;
   wire new_n9990_;
   wire new_n9989_;
   wire new_n9988_1_;
   wire new_n9987_;
   wire new_n9986_;
   wire new_n9985_1_;
   wire new_n9984_;
   wire new_n9983_;
   wire new_n9982_;
   wire new_n9981_1_;
   wire new_n9976_1_;
   wire new_n9975_;
   wire new_n9974_;
   wire new_n9973_;
   wire new_n9972_;
   wire new_n9971_1_;
   wire new_n9970_;
   wire new_n9969_;
   wire new_n9968_;
   wire new_n9967_;
   wire new_n9966_1_;
   wire new_n9965_;
   wire new_n9964_;
   wire new_n9963_;
   wire new_n9951_;
   wire new_n9950_;
   wire new_n9949_1_;
   wire new_n9939_1_;
   wire new_n9938_;
   wire new_n9935_1_;
   wire new_n9934_;
   wire new_n9933_;
   wire new_n9928_;
   wire new_n9927_;
   wire new_n9920_;
   wire new_n9919_;
   wire new_n9918_1_;
   wire new_n9917_;
   wire new_n9916_;
   wire new_n9915_;
   wire new_n9914_1_;
   wire new_n9910_;
   wire new_n9909_;
   wire new_n9908_;
   wire new_n9903_;
   wire new_n9902_1_;
   wire new_n9901_;
   wire new_n9900_;
   wire new_n9885_1_;
   wire new_n9883_;
   wire new_n9881_;
   wire new_n9876_;
   wire new_n9875_1_;
   wire new_n9874_;
   wire new_n9873_;
   wire new_n9872_;
   wire new_n9871_1_;
   wire new_n9870_;
   wire new_n9869_;
   wire new_n9868_;
   wire new_n9867_1_;
   wire new_n9866_;
   wire new_n9865_;
   wire new_n9857_;
   wire new_n9856_;
   wire new_n9855_;
   wire new_n9854_;
   wire new_n9853_1_;
   wire new_n9852_;
   wire new_n9851_;
   wire new_n9850_;
   wire new_n9849_1_;
   wire new_n9848_;
   wire new_n9847_;
   wire new_n9846_;
   wire new_n9844_1_;
   wire new_n9839_;
   wire new_n9838_;
   wire new_n9835_;
   wire new_n9834_;
   wire new_n9832_;
   wire new_n9831_;
   wire new_n9830_;
   wire new_n9829_;
   wire new_n9828_1_;
   wire new_n9826_;
   wire new_n9825_;
   wire new_n9822_;
   wire new_n9821_;
   wire new_n9813_;
   wire new_n9812_;
   wire new_n9810_;
   wire new_n9805_1_;
   wire new_n9804_;
   wire new_n9803_;
   wire new_n9798_;
   wire new_n9797_;
   wire new_n9794_;
   wire new_n9793_;
   wire new_n9791_;
   wire new_n9790_;
   wire new_n9789_;
   wire new_n9788_;
   wire new_n9787_1_;
   wire new_n9786_;
   wire new_n9785_;
   wire new_n9784_;
   wire new_n9783_1_;
   wire new_n9782_;
   wire new_n9781_;
   wire new_n9780_;
   wire new_n9779_;
   wire new_n9778_1_;
   wire new_n9777_;
   wire new_n9776_;
   wire new_n9775_;
   wire new_n9774_;
   wire new_n9773_1_;
   wire new_n9768_1_;
   wire new_n9767_;
   wire new_n9765_;
   wire new_n9764_;
   wire new_n9763_1_;
   wire new_n9762_;
   wire new_n9761_;
   wire new_n9760_;
   wire new_n9759_;
   wire new_n9758_1_;
   wire new_n9757_;
   wire new_n9755_;
   wire new_n9752_;
   wire new_n9747_;
   wire new_n9746_1_;
   wire new_n9745_;
   wire new_n9744_;
   wire new_n9743_;
   wire new_n9742_1_;
   wire new_n9741_;
   wire new_n9736_;
   wire new_n9735_;
   wire new_n9732_;
   wire new_n9731_;
   wire new_n9730_;
   wire new_n9729_1_;
   wire new_n9724_1_;
   wire new_n9723_;
   wire new_n9722_;
   wire new_n9721_;
   wire new_n9720_;
   wire new_n9718_;
   wire new_n9717_;
   wire new_n9708_;
   wire new_n9707_;
   wire new_n9703_;
   wire new_n9702_;
   wire new_n9694_;
   wire new_n9693_;
   wire new_n9686_;
   wire new_n9685_;
   wire new_n9684_;
   wire new_n9683_1_;
   wire new_n9682_;
   wire new_n9679_;
   wire new_n9678_1_;
   wire new_n9677_;
   wire new_n9676_;
   wire new_n9675_;
   wire new_n9674_;
   wire new_n9673_1_;
   wire new_n9670_;
   wire new_n9669_;
   wire new_n9668_1_;
   wire new_n9667_;
   wire new_n9666_;
   wire new_n9665_;
   wire new_n9664_1_;
   wire new_n9662_;
   wire new_n9661_;
   wire new_n9659_;
   wire new_n9651_1_;
   wire new_n9650_;
   wire new_n9649_;
   wire new_n9648_;
   wire new_n9647_1_;
   wire new_n9646_;
   wire new_n9645_;
   wire new_n9644_;
   wire new_n9643_;
   wire new_n9637_;
   wire new_n9636_;
   wire new_n9635_;
   wire new_n9634_;
   wire new_n9633_1_;
   wire new_n9632_;
   wire new_n9631_;
   wire new_n9630_;
   wire new_n9629_;
   wire new_n9628_1_;
   wire new_n9627_;
   wire new_n9623_;
   wire new_n9620_1_;
   wire new_n9619_;
   wire new_n9618_;
   wire new_n9613_;
   wire new_n9612_;
   wire new_n9611_1_;
   wire new_n9610_;
   wire new_n9608_;
   wire new_n9607_;
   wire new_n9604_;
   wire new_n9602_1_;
   wire new_n9601_;
   wire new_n9594_;
   wire new_n9593_;
   wire new_n9591_;
   wire new_n9590_;
   wire new_n9587_;
   wire new_n9586_;
   wire new_n9584_;
   wire new_n9583_1_;
   wire new_n9581_;
   wire new_n9580_;
   wire new_n9574_1_;
   wire new_n9573_;
   wire new_n9571_;
   wire new_n9570_;
   wire new_n9569_1_;
   wire new_n9562_;
   wire new_n9561_;
   wire new_n9560_;
   wire new_n9559_1_;
   wire new_n9558_;
   wire new_n9546_1_;
   wire new_n9541_1_;
   wire new_n9540_;
   wire new_n9539_;
   wire new_n9538_;
   wire new_n9537_1_;
   wire new_n9536_;
   wire new_n9531_;
   wire new_n9530_;
   wire new_n9529_;
   wire new_n9528_1_;
   wire new_n9527_;
   wire new_n9526_;
   wire new_n9525_1_;
   wire new_n9524_;
   wire new_n9523_;
   wire new_n9522_;
   wire new_n9520_1_;
   wire new_n9517_1_;
   wire new_n9516_;
   wire new_n9509_;
   wire new_n9508_;
   wire new_n9507_1_;
   wire new_n9504_;
   wire new_n9503_;
   wire new_n9502_1_;
   wire new_n9501_;
   wire new_n9498_;
   wire new_n9497_1_;
   wire new_n9496_;
   wire new_n9495_;
   wire new_n9494_;
   wire new_n9493_;
   wire new_n9492_1_;
   wire new_n9491_;
   wire new_n9490_;
   wire new_n9489_;
   wire new_n9488_;
   wire new_n9487_1_;
   wire new_n9486_;
   wire new_n9485_;
   wire new_n9484_;
   wire new_n9481_;
   wire new_n9480_;
   wire new_n9478_1_;
   wire new_n9477_;
   wire new_n9469_;
   wire new_n9468_;
   wire new_n9467_1_;
   wire new_n9465_;
   wire new_n9464_;
   wire new_n9463_;
   wire new_n9462_1_;
   wire new_n9458_;
   wire new_n9457_;
   wire new_n9453_;
   wire new_n9452_;
   wire new_n9451_;
   wire new_n9450_;
   wire new_n9449_1_;
   wire new_n9448_;
   wire new_n9447_;
   wire new_n9446_;
   wire new_n9445_1_;
   wire new_n9442_;
   wire new_n9441_1_;
   wire new_n9440_;
   wire new_n9439_;
   wire new_n9438_;
   wire new_n9436_1_;
   wire new_n9435_;
   wire new_n9434_;
   wire new_n9433_;
   wire new_n9428_1_;
   wire new_n9427_;
   wire new_n9426_;
   wire new_n9421_;
   wire new_n9420_1_;
   wire new_n9417_;
   wire new_n9416_;
   wire new_n9405_1_;
   wire new_n9404_;
   wire new_n9403_;
   wire new_n9401_;
   wire new_n9400_;
   wire new_n9393_1_;
   wire new_n9392_;
   wire new_n9391_;
   wire new_n9387_;
   wire new_n9385_1_;
   wire new_n9384_;
   wire new_n9381_1_;
   wire new_n9380_;
   wire new_n9378_;
   wire new_n9377_1_;
   wire new_n9376_;
   wire new_n9375_;
   wire new_n9374_;
   wire new_n9371_;
   wire new_n9370_1_;
   wire new_n9367_;
   wire new_n9366_;
   wire new_n9360_;
   wire new_n9359_;
   wire new_n9358_;
   wire new_n9357_;
   wire new_n9356_1_;
   wire new_n9355_;
   wire new_n9354_;
   wire new_n9351_;
   wire new_n9349_;
   wire new_n9348_1_;
   wire new_n9347_;
   wire new_n9345_;
   wire new_n9344_;
   wire new_n9343_1_;
   wire new_n9342_;
   wire new_n9341_;
   wire new_n9340_;
   wire new_n9339_1_;
   wire new_n9338_;
   wire new_n9333_;
   wire new_n9332_;
   wire new_n9331_;
   wire new_n9330_1_;
   wire new_n9329_;
   wire new_n9328_;
   wire new_n9327_;
   wire new_n9326_1_;
   wire new_n9325_;
   wire new_n9324_;
   wire new_n9323_;
   wire new_n9322_;
   wire new_n9321_1_;
   wire new_n9320_;
   wire new_n9316_1_;
   wire new_n9315_;
   wire new_n9311_;
   wire new_n9310_;
   wire new_n9308_;
   wire new_n9307_1_;
   wire new_n9306_;
   wire new_n9305_;
   wire new_n9304_;
   wire new_n9303_;
   wire new_n9289_;
   wire new_n9288_;
   wire new_n9285_;
   wire new_n9284_;
   wire new_n9283_;
   wire new_n9282_1_;
   wire new_n9281_;
   wire new_n9280_;
   wire new_n9279_;
   wire new_n9278_;
   wire new_n9277_1_;
   wire new_n9276_;
   wire new_n9275_;
   wire new_n9274_;
   wire new_n9273_;
   wire new_n9272_1_;
   wire new_n9271_;
   wire new_n9270_;
   wire new_n9269_;
   wire new_n9268_;
   wire new_n9267_1_;
   wire new_n9262_;
   wire new_n9261_;
   wire new_n9257_;
   wire new_n9256_;
   wire new_n9255_;
   wire new_n9254_1_;
   wire new_n9253_;
   wire new_n9252_;
   wire new_n9251_;
   wire new_n9250_1_;
   wire new_n9249_;
   wire new_n9248_;
   wire new_n9247_;
   wire new_n9243_;
   wire new_n9242_1_;
   wire new_n9241_;
   wire new_n9240_;
   wire new_n9239_;
   wire new_n9238_1_;
   wire new_n9237_;
   wire new_n9236_;
   wire new_n9235_;
   wire new_n9234_;
   wire new_n9233_1_;
   wire new_n9232_;
   wire new_n9231_;
   wire new_n9230_;
   wire new_n9228_1_;
   wire new_n9227_;
   wire new_n9226_;
   wire new_n9225_1_;
   wire new_n9224_;
   wire new_n9223_;
   wire new_n9222_;
   wire new_n9221_;
   wire new_n9220_1_;
   wire new_n9219_;
   wire new_n9218_;
   wire new_n9217_;
   wire new_n9216_;
   wire new_n9215_1_;
   wire new_n9211_1_;
   wire new_n9210_;
   wire new_n9205_;
   wire new_n9204_;
   wire new_n9203_;
   wire new_n9197_;
   wire new_n9196_1_;
   wire new_n9195_;
   wire new_n9193_;
   wire new_n9192_1_;
   wire new_n9191_;
   wire new_n9190_;
   wire new_n9189_;
   wire new_n9188_;
   wire new_n9187_1_;
   wire new_n9186_;
   wire new_n9185_;
   wire new_n9184_;
   wire new_n9183_;
   wire new_n9182_1_;
   wire new_n9181_;
   wire new_n9180_;
   wire new_n9179_;
   wire new_n9178_1_;
   wire new_n9177_;
   wire new_n9176_;
   wire new_n9175_;
   wire new_n9174_;
   wire new_n9173_1_;
   wire new_n9172_;
   wire new_n9171_;
   wire new_n9170_;
   wire new_n9163_;
   wire new_n9162_;
   wire new_n9161_;
   wire new_n9160_1_;
   wire new_n9159_;
   wire new_n9158_;
   wire new_n9156_1_;
   wire new_n9155_;
   wire new_n9149_;
   wire new_n9148_;
   wire new_n9147_;
   wire new_n9146_1_;
   wire new_n9145_;
   wire new_n9144_;
   wire new_n9143_1_;
   wire new_n9142_;
   wire new_n9141_;
   wire new_n9140_;
   wire new_n9139_;
   wire new_n9138_1_;
   wire new_n9137_;
   wire new_n9136_;
   wire new_n9135_;
   wire new_n9127_;
   wire new_n9126_;
   wire new_n9125_;
   wire new_n9124_1_;
   wire new_n9123_;
   wire new_n9122_;
   wire new_n9121_;
   wire new_n9120_1_;
   wire new_n9119_;
   wire new_n9118_;
   wire new_n9117_;
   wire new_n9116_;
   wire new_n9113_;
   wire new_n9112_;
   wire new_n9111_;
   wire new_n9110_1_;
   wire new_n9109_;
   wire new_n9108_;
   wire new_n9107_;
   wire new_n9106_1_;
   wire new_n9105_;
   wire new_n9103_;
   wire new_n9102_;
   wire new_n9098_;
   wire new_n9097_;
   wire new_n9096_1_;
   wire new_n9095_;
   wire new_n9094_;
   wire new_n9093_;
   wire new_n9092_;
   wire new_n9091_1_;
   wire new_n9090_;
   wire new_n9089_;
   wire new_n9088_;
   wire new_n9087_;
   wire new_n9086_1_;
   wire new_n9085_;
   wire new_n9084_;
   wire new_n9083_;
   wire new_n9082_1_;
   wire new_n9081_;
   wire new_n9080_;
   wire new_n9073_;
   wire new_n9072_;
   wire new_n9071_;
   wire new_n9070_;
   wire new_n9069_1_;
   wire new_n9068_;
   wire new_n9067_;
   wire new_n9066_;
   wire new_n9065_1_;
   wire new_n9058_;
   wire new_n9057_1_;
   wire new_n9056_;
   wire new_n9055_;
   wire new_n9054_;
   wire new_n9053_;
   wire new_n9052_1_;
   wire new_n9051_;
   wire new_n9050_;
   wire new_n9049_;
   wire new_n9048_;
   wire new_n9047_1_;
   wire new_n9046_;
   wire new_n9045_;
   wire new_n9042_1_;
   wire new_n9039_;
   wire new_n9038_;
   wire new_n9037_1_;
   wire new_n9036_;
   wire new_n9035_;
   wire new_n9033_;
   wire new_n9032_;
   wire new_n9031_;
   wire new_n9030_1_;
   wire new_n9029_;
   wire new_n9028_;
   wire new_n9027_;
   wire new_n9026_;
   wire new_n9025_1_;
   wire new_n9024_;
   wire new_n9023_;
   wire new_n9022_1_;
   wire new_n9021_;
   wire new_n9020_;
   wire new_n9018_;
   wire new_n9017_1_;
   wire new_n9014_1_;
   wire new_n9013_;
   wire new_n9012_;
   wire new_n9009_;
   wire new_n9008_;
   wire new_n9003_;
   wire new_n9002_;
   wire new_n9001_;
   wire new_n8997_;
   wire new_n8996_;
   wire new_n8991_;
   wire new_n8990_1_;
   wire new_n8985_;
   wire new_n8984_;
   wire new_n8973_;
   wire new_n8972_;
   wire new_n8969_;
   wire new_n8968_;
   wire new_n8964_;
   wire new_n8963_1_;
   wire new_n8962_;
   wire new_n8959_;
   wire new_n8958_1_;
   wire new_n8957_;
   wire new_n8948_1_;
   wire new_n8947_;
   wire new_n8945_;
   wire new_n8944_;
   wire new_n8940_;
   wire new_n8939_1_;
   wire new_n8938_;
   wire new_n8937_;
   wire new_n8936_;
   wire new_n8935_;
   wire new_n8934_1_;
   wire new_n8933_;
   wire new_n8932_;
   wire new_n8931_1_;
   wire new_n8930_;
   wire new_n8929_;
   wire new_n8928_;
   wire new_n8927_;
   wire new_n8925_;
   wire new_n8924_;
   wire new_n8923_;
   wire new_n8922_1_;
   wire new_n8921_;
   wire new_n8920_;
   wire new_n8919_;
   wire new_n8916_;
   wire new_n8915_;
   wire new_n8913_;
   wire new_n8912_1_;
   wire new_n8911_;
   wire new_n8909_;
   wire new_n8908_1_;
   wire new_n8907_;
   wire new_n8905_;
   wire new_n8899_1_;
   wire new_n8898_;
   wire new_n8897_;
   wire new_n8888_;
   wire new_n8887_;
   wire new_n8886_1_;
   wire new_n8885_;
   wire new_n8884_;
   wire new_n8883_;
   wire new_n8882_1_;
   wire new_n8881_;
   wire new_n8880_;
   wire new_n8879_;
   wire new_n8878_;
   wire new_n8873_1_;
   wire new_n8872_;
   wire new_n8861_;
   wire new_n8860_1_;
   wire new_n8859_;
   wire new_n8858_;
   wire new_n8857_;
   wire new_n8854_;
   wire new_n8853_;
   wire new_n8852_;
   wire new_n8851_;
   wire new_n8848_;
   wire new_n8846_;
   wire new_n8845_1_;
   wire new_n8844_;
   wire new_n8843_;
   wire new_n8842_;
   wire new_n8841_;
   wire new_n8840_1_;
   wire new_n8839_;
   wire new_n8838_;
   wire new_n8837_;
   wire new_n8836_;
   wire new_n8835_1_;
   wire new_n8834_;
   wire new_n8833_;
   wire new_n8832_;
   wire new_n8831_1_;
   wire new_n8830_;
   wire new_n8829_;
   wire new_n8828_;
   wire new_n8822_;
   wire new_n8821_;
   wire new_n8817_;
   wire new_n8816_;
   wire new_n8810_;
   wire new_n8805_1_;
   wire new_n8804_;
   wire new_n8803_;
   wire new_n8802_;
   wire new_n8801_;
   wire new_n8800_1_;
   wire new_n8799_;
   wire new_n8798_;
   wire new_n8797_1_;
   wire new_n8796_;
   wire new_n8795_;
   wire new_n8794_;
   wire new_n8793_1_;
   wire new_n8792_;
   wire new_n8790_;
   wire new_n8789_;
   wire new_n8788_1_;
   wire new_n8782_;
   wire new_n8781_;
   wire new_n8780_1_;
   wire new_n8779_;
   wire new_n8778_;
   wire new_n8774_;
   wire new_n8773_;
   wire new_n8767_1_;
   wire new_n8766_;
   wire new_n8765_;
   wire new_n8764_;
   wire new_n8761_;
   wire new_n8760_;
   wire new_n8759_;
   wire new_n8758_;
   wire new_n8757_1_;
   wire new_n8756_;
   wire new_n8755_;
   wire new_n8754_;
   wire new_n8753_1_;
   wire new_n8747_;
   wire new_n8746_;
   wire new_n8745_;
   wire new_n8744_;
   wire new_n8743_1_;
   wire new_n8742_;
   wire new_n8741_;
   wire new_n8740_;
   wire new_n8739_1_;
   wire new_n8738_;
   wire new_n8737_;
   wire new_n8736_;
   wire new_n8735_;
   wire new_n8734_1_;
   wire new_n8733_;
   wire new_n8732_;
   wire new_n8731_;
   wire new_n8730_1_;
   wire new_n8729_;
   wire new_n8728_;
   wire new_n8727_;
   wire new_n8726_;
   wire new_n8725_1_;
   wire new_n8724_;
   wire new_n8723_;
   wire new_n8719_;
   wire new_n8718_;
   wire new_n8717_;
   wire new_n8713_;
   wire new_n8712_;
   wire new_n8700_;
   wire new_n8698_1_;
   wire new_n8696_;
   wire new_n8695_;
   wire new_n8694_1_;
   wire new_n8692_;
   wire new_n8691_;
   wire new_n8690_;
   wire new_n8687_;
   wire new_n8686_;
   wire new_n8685_1_;
   wire new_n8681_1_;
   wire new_n8680_;
   wire new_n8679_;
   wire new_n8678_;
   wire new_n8677_;
   wire new_n8675_;
   wire new_n8671_1_;
   wire new_n8670_;
   wire new_n8669_;
   wire new_n8668_;
   wire new_n8667_;
   wire new_n8666_1_;
   wire new_n8665_;
   wire new_n8664_;
   wire new_n8663_;
   wire new_n8662_1_;
   wire new_n8661_;
   wire new_n8660_;
   wire new_n8659_;
   wire new_n8658_1_;
   wire new_n8657_;
   wire new_n8656_;
   wire new_n8655_;
   wire new_n8654_1_;
   wire new_n8653_;
   wire new_n8652_;
   wire new_n8651_;
   wire new_n8650_1_;
   wire new_n8649_;
   wire new_n8648_;
   wire new_n8646_;
   wire new_n8645_1_;
   wire new_n8643_;
   wire new_n8642_;
   wire new_n8641_1_;
   wire new_n8637_1_;
   wire new_n8636_;
   wire new_n8629_;
   wire new_n8628_1_;
   wire new_n8626_;
   wire new_n8625_1_;
   wire new_n8622_;
   wire new_n8621_1_;
   wire new_n8620_;
   wire new_n8619_;
   wire new_n8618_;
   wire new_n8617_;
   wire new_n8616_1_;
   wire new_n8615_;
   wire new_n8614_;
   wire new_n8613_;
   wire new_n8612_1_;
   wire new_n8611_;
   wire new_n8610_;
   wire new_n8609_;
   wire new_n8608_;
   wire new_n8601_;
   wire new_n8600_;
   wire new_n8599_;
   wire new_n8598_1_;
   wire new_n8597_;
   wire new_n8596_;
   wire new_n8594_;
   wire new_n8593_1_;
   wire new_n8592_;
   wire new_n8591_;
   wire new_n8587_;
   wire new_n8586_;
   wire new_n8581_;
   wire new_n8580_;
   wire new_n8579_;
   wire new_n8578_1_;
   wire new_n8577_;
   wire new_n8576_;
   wire new_n8575_1_;
   wire new_n8574_;
   wire new_n8573_;
   wire new_n8572_;
   wire new_n8571_;
   wire new_n8570_1_;
   wire new_n8569_;
   wire new_n8568_;
   wire new_n8566_;
   wire new_n8565_1_;
   wire new_n8561_1_;
   wire new_n8560_;
   wire new_n8559_;
   wire new_n8556_;
   wire new_n8555_;
   wire new_n8554_;
   wire new_n8553_;
   wire new_n8552_1_;
   wire new_n8551_;
   wire new_n8550_;
   wire new_n8549_1_;
   wire new_n8548_;
   wire new_n8547_;
   wire new_n8546_;
   wire new_n8545_;
   wire new_n8543_;
   wire new_n8541_;
   wire new_n8540_1_;
   wire new_n8536_;
   wire new_n8535_1_;
   wire new_n8534_;
   wire new_n8533_;
   wire new_n8532_;
   wire new_n8531_1_;
   wire new_n8530_;
   wire new_n8529_;
   wire new_n8528_;
   wire new_n8527_;
   wire new_n8526_1_;
   wire new_n8525_;
   wire new_n8524_;
   wire new_n8523_;
   wire new_n8522_1_;
   wire new_n8521_;
   wire new_n8520_;
   wire new_n8519_;
   wire new_n8518_;
   wire new_n8517_1_;
   wire new_n8516_;
   wire new_n8515_;
   wire new_n8514_;
   wire new_n8513_1_;
   wire new_n8505_;
   wire new_n8503_;
   wire new_n8502_;
   wire new_n8501_;
   wire new_n8500_;
   wire new_n8499_1_;
   wire new_n8498_;
   wire new_n8497_;
   wire new_n8496_;
   wire new_n8495_;
   wire new_n8494_1_;
   wire new_n8493_;
   wire new_n8492_;
   wire new_n8491_1_;
   wire new_n8490_;
   wire new_n8489_;
   wire new_n8488_;
   wire new_n8487_;
   wire new_n8486_1_;
   wire new_n8485_;
   wire new_n8484_;
   wire new_n8483_;
   wire new_n8482_;
   wire new_n8481_1_;
   wire new_n8480_;
   wire new_n8475_;
   wire new_n8474_;
   wire new_n8473_;
   wire new_n8469_;
   wire new_n8468_;
   wire new_n8463_;
   wire new_n8461_;
   wire new_n8460_;
   wire new_n8459_1_;
   wire new_n8458_;
   wire new_n8457_;
   wire new_n8456_;
   wire new_n8455_1_;
   wire new_n8454_;
   wire new_n8453_;
   wire new_n8452_;
   wire new_n8451_1_;
   wire new_n8450_;
   wire new_n8449_;
   wire new_n8448_;
   wire new_n8447_1_;
   wire new_n8446_;
   wire new_n8445_;
   wire new_n8444_;
   wire new_n8443_1_;
   wire new_n8441_;
   wire new_n8440_;
   wire new_n8439_;
   wire new_n8438_1_;
   wire new_n8436_;
   wire new_n8435_1_;
   wire new_n8431_;
   wire new_n8430_1_;
   wire new_n8429_;
   wire new_n8428_;
   wire new_n8427_;
   wire new_n8426_1_;
   wire new_n8425_;
   wire new_n8424_;
   wire new_n8423_;
   wire new_n8422_1_;
   wire new_n8421_;
   wire new_n8420_;
   wire new_n8419_;
   wire new_n8418_1_;
   wire new_n8416_;
   wire new_n8415_1_;
   wire new_n8412_;
   wire new_n8411_;
   wire new_n8410_1_;
   wire new_n8407_;
   wire new_n8406_;
   wire new_n8405_1_;
   wire new_n8404_;
   wire new_n8403_;
   wire new_n8402_;
   wire new_n8401_1_;
   wire new_n8400_;
   wire new_n8396_1_;
   wire new_n8395_;
   wire new_n8394_;
   wire new_n8393_;
   wire new_n8392_1_;
   wire new_n8391_;
   wire new_n8390_;
   wire new_n8389_;
   wire new_n8387_1_;
   wire new_n8386_;
   wire new_n8383_;
   wire new_n8382_1_;
   wire new_n8381_;
   wire new_n8380_;
   wire new_n8379_;
   wire new_n8377_1_;
   wire new_n8376_;
   wire new_n8375_;
   wire new_n8374_;
   wire new_n8373_;
   wire new_n8372_1_;
   wire new_n8371_;
   wire new_n8370_;
   wire new_n8369_;
   wire new_n8368_;
   wire new_n8367_1_;
   wire new_n8366_;
   wire new_n8365_;
   wire new_n8364_;
   wire new_n8363_;
   wire new_n8362_1_;
   wire new_n8361_;
   wire new_n8360_;
   wire new_n8359_1_;
   wire new_n8358_;
   wire new_n8357_;
   wire new_n8356_;
   wire new_n8355_;
   wire new_n8354_1_;
   wire new_n8350_1_;
   wire new_n8349_;
   wire new_n8348_;
   wire new_n8347_;
   wire new_n8346_;
   wire new_n8345_1_;
   wire new_n8344_;
   wire new_n8343_;
   wire new_n8342_;
   wire new_n8341_;
   wire new_n8339_;
   wire new_n8338_;
   wire new_n8336_;
   wire new_n8335_;
   wire new_n8334_1_;
   wire new_n8327_;
   wire new_n8326_;
   wire new_n8325_;
   wire new_n8324_1_;
   wire new_n8307_1_;
   wire new_n8306_;
   wire new_n8305_;
   wire new_n8304_;
   wire new_n8303_1_;
   wire new_n8301_;
   wire new_n8300_;
   wire new_n8299_1_;
   wire new_n8298_;
   wire new_n8297_;
   wire new_n8296_;
   wire new_n8294_1_;
   wire new_n8293_;
   wire new_n8292_;
   wire new_n8291_;
   wire new_n8289_1_;
   wire new_n8288_;
   wire new_n8285_;
   wire new_n8284_1_;
   wire new_n8282_;
   wire new_n8281_;
   wire new_n8280_1_;
   wire new_n8276_1_;
   wire new_n8275_;
   wire new_n8274_;
   wire new_n8273_;
   wire new_n8272_;
   wire new_n8271_1_;
   wire new_n8270_;
   wire new_n8269_;
   wire new_n8267_;
   wire new_n8266_1_;
   wire new_n8265_;
   wire new_n8263_;
   wire new_n8262_1_;
   wire new_n8254_;
   wire new_n8253_1_;
   wire new_n8252_;
   wire new_n8251_;
   wire new_n8250_;
   wire new_n8249_1_;
   wire new_n8248_;
   wire new_n8247_;
   wire new_n8246_;
   wire new_n8245_1_;
   wire new_n8244_;
   wire new_n8243_;
   wire new_n8234_;
   wire new_n8233_;
   wire new_n8231_;
   wire new_n8230_;
   wire new_n8229_;
   wire new_n8228_1_;
   wire new_n8225_;
   wire new_n8224_1_;
   wire new_n8221_;
   wire new_n8220_1_;
   wire new_n8219_;
   wire new_n8218_;
   wire new_n8217_;
   wire new_n8216_1_;
   wire new_n8215_;
   wire new_n8214_;
   wire new_n8212_;
   wire new_n8211_1_;
   wire new_n8210_;
   wire new_n8209_;
   wire new_n8208_;
   wire new_n8207_;
   wire new_n8206_1_;
   wire new_n8205_;
   wire new_n8204_;
   wire new_n8203_;
   wire new_n8202_1_;
   wire new_n8201_;
   wire new_n8200_;
   wire new_n8199_;
   wire new_n8198_;
   wire new_n8197_1_;
   wire new_n8193_;
   wire new_n8192_1_;
   wire new_n8191_;
   wire new_n8188_1_;
   wire new_n8187_;
   wire new_n8186_;
   wire new_n8185_;
   wire new_n8184_;
   wire new_n8183_1_;
   wire new_n8181_;
   wire new_n8180_;
   wire new_n8179_1_;
   wire new_n8178_;
   wire new_n8177_;
   wire new_n8176_;
   wire new_n8175_;
   wire new_n8174_1_;
   wire new_n8173_;
   wire new_n8172_;
   wire new_n8171_;
   wire new_n8170_1_;
   wire new_n8169_;
   wire new_n8168_;
   wire new_n8167_;
   wire new_n8166_1_;
   wire new_n8165_;
   wire new_n8164_;
   wire new_n8163_;
   wire new_n8162_;
   wire new_n8161_1_;
   wire new_n8160_;
   wire new_n8159_;
   wire new_n8158_;
   wire new_n8157_;
   wire new_n8156_1_;
   wire new_n8155_;
   wire new_n8154_;
   wire new_n8153_;
   wire new_n8151_;
   wire new_n8150_;
   wire new_n8149_;
   wire new_n8147_1_;
   wire new_n8146_;
   wire new_n8145_;
   wire new_n8144_1_;
   wire new_n8143_;
   wire new_n8142_;
   wire new_n8141_;
   wire new_n8140_1_;
   wire new_n8139_;
   wire new_n8135_1_;
   wire new_n8134_;
   wire new_n8133_;
   wire new_n8132_;
   wire new_n8131_;
   wire new_n8124_;
   wire new_n8123_;
   wire new_n8122_;
   wire new_n8121_1_;
   wire new_n8120_;
   wire new_n8119_;
   wire new_n8118_;
   wire new_n8117_;
   wire new_n8114_;
   wire new_n8113_;
   wire new_n8112_1_;
   wire new_n8107_1_;
   wire new_n8106_;
   wire new_n8105_;
   wire new_n8104_;
   wire new_n8103_;
   wire new_n8102_1_;
   wire new_n8100_;
   wire new_n8099_;
   wire new_n8091_;
   wire new_n8090_;
   wire new_n8084_;
   wire new_n8083_;
   wire new_n8082_;
   wire new_n8081_;
   wire new_n8080_1_;
   wire new_n8079_;
   wire new_n8078_;
   wire new_n8077_;
   wire new_n8076_;
   wire new_n8075_1_;
   wire new_n8074_;
   wire new_n8073_;
   wire new_n8072_1_;
   wire new_n8071_;
   wire new_n8068_;
   wire new_n8067_1_;
   wire new_n8066_;
   wire new_n8065_;
   wire new_n8064_1_;
   wire new_n8061_;
   wire new_n8060_;
   wire new_n8059_1_;
   wire new_n8058_;
   wire new_n8057_;
   wire new_n8056_1_;
   wire new_n8055_;
   wire new_n8054_;
   wire new_n8053_;
   wire new_n8052_;
   wire new_n8051_1_;
   wire new_n8050_;
   wire new_n8049_;
   wire new_n8048_;
   wire new_n8044_;
   wire new_n8043_;
   wire new_n8042_1_;
   wire new_n8041_;
   wire new_n8040_;
   wire new_n8035_;
   wire new_n8034_;
   wire new_n8033_1_;
   wire new_n8032_;
   wire new_n8031_;
   wire new_n8030_;
   wire new_n8029_;
   wire new_n8028_1_;
   wire new_n8027_;
   wire new_n8026_;
   wire new_n8025_;
   wire new_n8024_1_;
   wire new_n8023_;
   wire new_n8022_;
   wire new_n8021_;
   wire new_n8020_;
   wire new_n8011_;
   wire new_n8010_1_;
   wire new_n8009_;
   wire new_n8005_1_;
   wire new_n8004_;
   wire new_n8001_;
   wire new_n8000_;
   wire new_n7999_;
   wire new_n7993_;
   wire new_n7992_;
   wire new_n7991_;
   wire new_n7990_;
   wire new_n7989_1_;
   wire new_n7987_;
   wire new_n7986_;
   wire new_n7985_1_;
   wire new_n7983_;
   wire new_n7978_;
   wire new_n7977_;
   wire new_n7976_;
   wire new_n7975_1_;
   wire new_n7972_;
   wire new_n7971_;
   wire new_n7970_1_;
   wire new_n7965_;
   wire new_n7964_;
   wire new_n7963_;
   wire new_n7962_1_;
   wire new_n7961_;
   wire new_n7960_;
   wire new_n7957_;
   wire new_n7956_;
   wire new_n7955_1_;
   wire new_n7954_;
   wire new_n7953_;
   wire new_n7952_;
   wire new_n7951_;
   wire new_n7950_1_;
   wire new_n7949_;
   wire new_n7946_;
   wire new_n7945_1_;
   wire new_n7944_;
   wire new_n7943_;
   wire new_n7942_1_;
   wire new_n7941_;
   wire new_n7940_;
   wire new_n7939_;
   wire new_n7938_;
   wire new_n7937_1_;
   wire new_n7936_;
   wire new_n7935_;
   wire new_n7934_;
   wire new_n7931_;
   wire new_n7930_;
   wire new_n7929_1_;
   wire new_n7925_;
   wire new_n7924_1_;
   wire new_n7923_;
   wire new_n7922_;
   wire new_n7921_;
   wire new_n7920_1_;
   wire new_n7919_;
   wire new_n7918_;
   wire new_n7917_;
   wire new_n7916_1_;
   wire new_n7915_;
   wire new_n7914_;
   wire new_n7913_;
   wire new_n7912_;
   wire new_n7911_1_;
   wire new_n7910_;
   wire new_n7909_;
   wire new_n7908_;
   wire new_n7907_;
   wire new_n7906_1_;
   wire new_n7905_;
   wire new_n7904_;
   wire new_n7903_;
   wire new_n7902_1_;
   wire new_n7896_;
   wire new_n7895_;
   wire new_n7892_;
   wire new_n7891_;
   wire new_n7878_1_;
   wire new_n7876_;
   wire new_n7875_1_;
   wire new_n7874_;
   wire new_n7873_;
   wire new_n7872_;
   wire new_n7869_;
   wire new_n7868_;
   wire new_n7865_;
   wire new_n7864_;
   wire new_n7863_1_;
   wire new_n7862_;
   wire new_n7861_;
   wire new_n7860_;
   wire new_n7859_;
   wire new_n7858_1_;
   wire new_n7857_;
   wire new_n7856_;
   wire new_n7855_;
   wire new_n7854_;
   wire new_n7853_1_;
   wire new_n7851_;
   wire new_n7850_;
   wire new_n7849_;
   wire new_n7848_1_;
   wire new_n7847_;
   wire new_n7845_1_;
   wire new_n7844_;
   wire new_n7843_;
   wire new_n7842_;
   wire new_n7841_;
   wire new_n7840_1_;
   wire new_n7839_;
   wire new_n7838_;
   wire new_n7837_;
   wire new_n7836_;
   wire new_n7835_1_;
   wire new_n7834_;
   wire new_n7833_;
   wire new_n7832_;
   wire new_n7831_1_;
   wire new_n7830_;
   wire new_n7829_;
   wire new_n7828_;
   wire new_n7827_;
   wire new_n7826_1_;
   wire new_n7825_;
   wire new_n7824_;
   wire new_n7823_;
   wire new_n7822_1_;
   wire new_n7821_;
   wire new_n7820_;
   wire new_n7819_;
   wire new_n7818_1_;
   wire new_n7817_;
   wire new_n7816_;
   wire new_n7815_1_;
   wire new_n7814_;
   wire new_n7813_;
   wire new_n7812_;
   wire new_n7811_;
   wire new_n7810_1_;
   wire new_n7806_1_;
   wire new_n7805_;
   wire new_n7804_;
   wire new_n7798_1_;
   wire new_n7797_;
   wire new_n7796_;
   wire new_n7795_;
   wire new_n7794_;
   wire new_n7792_;
   wire new_n7791_;
   wire new_n7779_1_;
   wire new_n7775_;
   wire new_n7774_;
   wire new_n7773_1_;
   wire new_n7772_;
   wire new_n7771_;
   wire new_n7767_;
   wire new_n7766_;
   wire new_n7762_;
   wire new_n7761_;
   wire new_n7760_1_;
   wire new_n7756_1_;
   wire new_n7755_;
   wire new_n7754_;
   wire new_n7753_;
   wire new_n7752_;
   wire new_n7747_;
   wire new_n7744_;
   wire new_n7741_1_;
   wire new_n7740_;
   wire new_n7739_;
   wire new_n7738_;
   wire new_n7736_;
   wire new_n7735_;
   wire new_n7734_;
   wire new_n7733_;
   wire new_n7732_1_;
   wire new_n7731_;
   wire new_n7730_;
   wire new_n7721_;
   wire new_n7720_;
   wire new_n7719_1_;
   wire new_n7718_;
   wire new_n7717_;
   wire new_n7716_;
   wire new_n7715_;
   wire new_n7714_1_;
   wire new_n7713_;
   wire new_n7712_;
   wire new_n7711_;
   wire new_n7710_;
   wire new_n7709_1_;
   wire new_n7708_;
   wire new_n7702_;
   wire new_n7701_;
   wire new_n7700_1_;
   wire new_n7699_;
   wire new_n7698_;
   wire new_n7697_;
   wire new_n7696_;
   wire new_n7695_1_;
   wire new_n7694_;
   wire new_n7693_;
   wire new_n7692_;
   wire new_n7691_1_;
   wire new_n7690_;
   wire new_n7689_;
   wire new_n7688_;
   wire new_n7687_;
   wire new_n7686_1_;
   wire new_n7685_;
   wire new_n7684_;
   wire new_n7683_;
   wire new_n7682_;
   wire new_n7681_1_;
   wire new_n7680_;
   wire new_n7679_;
   wire new_n7678_;
   wire new_n7677_;
   wire new_n7676_1_;
   wire new_n7675_;
   wire new_n7674_;
   wire new_n7669_;
   wire new_n7668_;
   wire new_n7667_;
   wire new_n7666_1_;
   wire new_n7665_;
   wire new_n7662_;
   wire new_n7661_1_;
   wire new_n7657_;
   wire new_n7656_;
   wire new_n7655_;
   wire new_n7652_;
   wire new_n7651_;
   wire new_n7650_;
   wire new_n7649_1_;
   wire new_n7648_;
   wire new_n7647_;
   wire new_n7646_;
   wire new_n7645_;
   wire new_n7644_1_;
   wire new_n7643_;
   wire new_n7633_;
   wire new_n7632_;
   wire new_n7631_1_;
   wire new_n7630_;
   wire new_n7629_;
   wire new_n7626_1_;
   wire new_n7625_;
   wire new_n7624_;
   wire new_n7623_;
   wire new_n7622_1_;
   wire new_n7621_;
   wire new_n7620_;
   wire new_n7619_;
   wire new_n7618_1_;
   wire new_n7617_;
   wire new_n7616_;
   wire new_n7615_;
   wire new_n7614_;
   wire new_n7613_1_;
   wire new_n7612_;
   wire new_n7609_;
   wire new_n7608_1_;
   wire new_n7605_;
   wire new_n7604_1_;
   wire new_n7602_;
   wire new_n7597_;
   wire new_n7596_1_;
   wire new_n7595_;
   wire new_n7594_;
   wire new_n7593_;
   wire new_n7590_;
   wire new_n7589_;
   wire new_n7588_;
   wire new_n7587_;
   wire new_n7586_1_;
   wire new_n7585_;
   wire new_n7584_;
   wire new_n7583_;
   wire new_n7582_;
   wire new_n7581_1_;
   wire new_n7580_;
   wire new_n7579_;
   wire new_n7578_;
   wire new_n7577_1_;
   wire new_n7576_;
   wire new_n7575_;
   wire new_n7574_;
   wire new_n7573_;
   wire new_n7572_1_;
   wire new_n7571_;
   wire new_n7570_;
   wire new_n7569_;
   wire new_n7568_;
   wire new_n7567_1_;
   wire new_n7566_;
   wire new_n7565_;
   wire new_n7564_;
   wire new_n7563_1_;
   wire new_n7562_;
   wire new_n7561_;
   wire new_n7560_;
   wire new_n7559_;
   wire new_n7558_1_;
   wire new_n7557_;
   wire new_n7556_;
   wire new_n7555_;
   wire new_n7554_;
   wire new_n7553_1_;
   wire new_n7552_;
   wire new_n7547_;
   wire new_n7545_;
   wire new_n7544_;
   wire new_n7543_1_;
   wire new_n7542_;
   wire new_n7541_;
   wire new_n7540_;
   wire new_n7538_;
   wire new_n7537_;
   wire new_n7533_;
   wire new_n7532_;
   wire new_n7531_;
   wire new_n7530_1_;
   wire new_n7529_;
   wire new_n7527_1_;
   wire new_n7526_;
   wire new_n7525_;
   wire new_n7523_;
   wire new_n7522_1_;
   wire new_n7521_;
   wire new_n7516_;
   wire new_n7515_;
   wire new_n7513_1_;
   wire new_n7512_;
   wire new_n7511_;
   wire new_n7510_;
   wire new_n7509_1_;
   wire new_n7508_;
   wire new_n7504_;
   wire new_n7503_;
   wire new_n7502_;
   wire new_n7501_1_;
   wire new_n7500_;
   wire new_n7499_;
   wire new_n7497_;
   wire new_n7496_1_;
   wire new_n7495_;
   wire new_n7494_;
   wire new_n7493_;
   wire new_n7492_1_;
   wire new_n7486_;
   wire new_n7485_;
   wire new_n7484_;
   wire new_n7483_;
   wire new_n7482_1_;
   wire new_n7472_;
   wire new_n7471_;
   wire new_n7467_;
   wire new_n7466_;
   wire new_n7465_;
   wire new_n7461_;
   wire new_n7460_;
   wire new_n7459_1_;
   wire new_n7452_;
   wire new_n7451_;
   wire new_n7450_1_;
   wire new_n7449_;
   wire new_n7448_;
   wire new_n7447_;
   wire new_n7446_1_;
   wire new_n7445_;
   wire new_n7444_;
   wire new_n7443_;
   wire new_n7442_1_;
   wire new_n7437_1_;
   wire new_n7436_;
   wire new_n7435_;
   wire new_n7430_;
   wire new_n7429_;
   wire new_n7428_;
   wire new_n7427_1_;
   wire new_n7424_;
   wire new_n7423_;
   wire new_n7422_1_;
   wire new_n7418_;
   wire new_n7417_1_;
   wire new_n7416_;
   wire new_n7415_;
   wire new_n7414_;
   wire new_n7413_1_;
   wire new_n7412_;
   wire new_n7411_;
   wire new_n7408_1_;
   wire new_n7407_;
   wire new_n7404_1_;
   wire new_n7403_;
   wire new_n7401_;
   wire new_n7400_1_;
   wire new_n7399_;
   wire new_n7398_;
   wire new_n7397_;
   wire new_n7396_;
   wire new_n7395_1_;
   wire new_n7394_;
   wire new_n7393_;
   wire new_n7392_;
   wire new_n7391_1_;
   wire new_n7390_;
   wire new_n7389_;
   wire new_n7388_;
   wire new_n7387_;
   wire new_n7386_1_;
   wire new_n7385_;
   wire new_n7384_;
   wire new_n7383_;
   wire new_n7382_;
   wire new_n7381_1_;
   wire new_n7380_;
   wire new_n7379_;
   wire new_n7378_;
   wire new_n7377_;
   wire new_n7376_1_;
   wire new_n7375_;
   wire new_n7374_;
   wire new_n7373_;
   wire new_n7372_1_;
   wire new_n7371_;
   wire new_n7370_;
   wire new_n7369_;
   wire new_n7368_1_;
   wire new_n7367_;
   wire new_n7366_;
   wire new_n7365_;
   wire new_n7364_;
   wire new_n7363_1_;
   wire new_n7362_;
   wire new_n7361_;
   wire new_n7360_;
   wire new_n7359_1_;
   wire new_n7358_;
   wire new_n7357_;
   wire new_n7356_;
   wire new_n7355_;
   wire new_n7354_1_;
   wire new_n7352_;
   wire new_n7351_;
   wire new_n7350_;
   wire new_n7346_;
   wire new_n7345_;
   wire new_n7344_1_;
   wire new_n7343_;
   wire new_n7342_;
   wire new_n7341_;
   wire new_n7340_1_;
   wire new_n7339_;
   wire new_n7337_;
   wire new_n7336_;
   wire new_n7335_1_;
   wire new_n7334_;
   wire new_n7333_;
   wire new_n7329_;
   wire new_n7328_;
   wire new_n7326_1_;
   wire new_n7325_;
   wire new_n7323_;
   wire new_n7322_;
   wire new_n7321_1_;
   wire new_n7320_;
   wire new_n7319_;
   wire new_n7312_1_;
   wire new_n7311_;
   wire new_n7310_;
   wire new_n7309_;
   wire new_n7306_;
   wire new_n7305_;
   wire new_n7304_;
   wire new_n7303_;
   wire new_n7302_1_;
   wire new_n7301_;
   wire new_n7300_;
   wire new_n7299_;
   wire new_n7298_;
   wire new_n7297_1_;
   wire new_n7296_;
   wire new_n7295_;
   wire new_n7294_;
   wire new_n7292_1_;
   wire new_n7291_;
   wire new_n7290_;
   wire new_n7289_;
   wire new_n7288_1_;
   wire new_n7287_;
   wire new_n7285_;
   wire new_n7284_1_;
   wire new_n7283_;
   wire new_n7282_;
   wire new_n7279_;
   wire new_n7278_;
   wire new_n7277_;
   wire new_n7276_;
   wire new_n7275_1_;
   wire new_n7274_;
   wire new_n7273_;
   wire new_n7272_;
   wire new_n7271_;
   wire new_n7270_1_;
   wire new_n7269_;
   wire new_n7268_;
   wire new_n7265_1_;
   wire new_n7264_;
   wire new_n7262_;
   wire new_n7258_;
   wire new_n7257_;
   wire new_n7256_1_;
   wire new_n7255_;
   wire new_n7254_;
   wire new_n7253_;
   wire new_n7252_1_;
   wire new_n7251_;
   wire new_n7250_;
   wire new_n7249_1_;
   wire new_n7248_;
   wire new_n7239_;
   wire new_n7236_;
   wire new_n7235_1_;
   wire new_n7234_;
   wire new_n7233_;
   wire new_n7232_;
   wire new_n7230_1_;
   wire new_n7229_;
   wire new_n7228_;
   wire new_n7227_;
   wire new_n7225_;
   wire new_n7224_;
   wire new_n7223_;
   wire new_n7222_;
   wire new_n7221_1_;
   wire new_n7220_;
   wire new_n7219_;
   wire new_n7218_;
   wire new_n7216_1_;
   wire new_n7215_;
   wire new_n7214_;
   wire new_n7213_;
   wire new_n7211_;
   wire new_n7210_;
   wire new_n7209_;
   wire new_n7208_;
   wire new_n7207_1_;
   wire new_n7206_;
   wire new_n7205_;
   wire new_n7204_;
   wire new_n7203_1_;
   wire new_n7202_;
   wire new_n7201_;
   wire new_n7200_;
   wire new_n7199_1_;
   wire new_n7198_;
   wire new_n7197_;
   wire new_n7196_;
   wire new_n7195_;
   wire new_n7194_1_;
   wire new_n7193_;
   wire new_n7192_;
   wire new_n7191_;
   wire new_n7190_1_;
   wire new_n7189_;
   wire new_n7188_;
   wire new_n7187_;
   wire new_n7186_;
   wire new_n7184_;
   wire new_n7183_;
   wire new_n7182_1_;
   wire new_n7181_;
   wire new_n7179_;
   wire new_n7178_;
   wire new_n7177_1_;
   wire new_n7175_;
   wire new_n7174_;
   wire new_n7173_;
   wire new_n7172_1_;
   wire new_n7171_;
   wire new_n7170_;
   wire new_n7169_;
   wire new_n7168_;
   wire new_n7167_1_;
   wire new_n7166_;
   wire new_n7165_;
   wire new_n7164_1_;
   wire new_n7163_;
   wire new_n7162_;
   wire new_n7161_;
   wire new_n7160_1_;
   wire new_n7159_;
   wire new_n7158_;
   wire new_n7157_;
   wire new_n7156_;
   wire new_n7155_1_;
   wire new_n7154_;
   wire new_n7153_;
   wire new_n7152_;
   wire new_n7151_1_;
   wire new_n7148_;
   wire new_n7137_;
   wire new_n7136_;
   wire new_n7135_;
   wire new_n7134_;
   wire new_n7133_1_;
   wire new_n7132_;
   wire new_n7131_;
   wire new_n7130_;
   wire new_n7129_;
   wire new_n7128_1_;
   wire new_n7127_;
   wire new_n7126_;
   wire new_n7125_1_;
   wire new_n7124_;
   wire new_n7123_;
   wire new_n7122_;
   wire new_n7121_;
   wire new_n7120_1_;
   wire new_n7119_;
   wire new_n7118_;
   wire new_n7117_;
   wire new_n7116_1_;
   wire new_n7115_;
   wire new_n7114_;
   wire new_n7113_;
   wire new_n7111_1_;
   wire new_n7110_;
   wire new_n7109_;
   wire new_n7108_;
   wire new_n7107_1_;
   wire new_n7106_;
   wire new_n7105_;
   wire new_n7104_;
   wire new_n7103_;
   wire new_n7102_1_;
   wire new_n7101_;
   wire new_n7100_;
   wire new_n7099_;
   wire new_n7098_1_;
   wire new_n7097_;
   wire new_n7093_1_;
   wire new_n7092_;
   wire new_n7091_;
   wire new_n7090_;
   wire new_n7089_1_;
   wire new_n7088_;
   wire new_n7087_;
   wire new_n7086_;
   wire new_n7085_1_;
   wire new_n7084_;
   wire new_n7083_;
   wire new_n7082_1_;
   wire new_n7081_;
   wire new_n7080_;
   wire new_n7079_;
   wire new_n7078_;
   wire new_n7077_1_;
   wire new_n7076_;
   wire new_n7075_;
   wire new_n7074_;
   wire new_n7073_;
   wire new_n7072_1_;
   wire new_n7071_;
   wire new_n7070_;
   wire new_n7069_;
   wire new_n7068_;
   wire new_n7067_1_;
   wire new_n7066_;
   wire new_n7065_;
   wire new_n7064_;
   wire new_n7063_;
   wire new_n7062_1_;
   wire new_n7061_;
   wire new_n7060_;
   wire new_n7059_;
   wire new_n7058_1_;
   wire new_n7057_;
   wire new_n7056_;
   wire new_n7055_;
   wire new_n7054_;
   wire new_n7053_1_;
   wire new_n7052_;
   wire new_n7051_;
   wire new_n7050_;
   wire new_n7049_1_;
   wire new_n7048_;
   wire new_n7047_;
   wire new_n7046_;
   wire new_n7045_1_;
   wire new_n7044_;
   wire new_n7043_;
   wire new_n7042_;
   wire new_n7035_;
   wire new_n7034_;
   wire new_n7029_;
   wire new_n7028_;
   wire new_n7027_1_;
   wire new_n7026_;
   wire new_n7025_;
   wire new_n7024_;
   wire new_n7023_1_;
   wire new_n7022_;
   wire new_n7021_;
   wire new_n7020_;
   wire new_n7019_;
   wire new_n7018_1_;
   wire new_n7017_;
   wire new_n7014_;
   wire new_n7013_1_;
   wire new_n7012_;
   wire new_n7011_;
   wire new_n7010_;
   wire new_n7009_1_;
   wire new_n7008_;
   wire new_n7007_;
   wire new_n7006_;
   wire new_n7005_1_;
   wire new_n7004_;
   wire new_n7003_;
   wire new_n7002_;
   wire new_n7001_;
   wire new_n7000_1_;
   wire new_n6999_;
   wire new_n6998_;
   wire new_n6997_;
   wire new_n6996_;
   wire new_n6995_1_;
   wire new_n6994_;
   wire new_n6993_;
   wire new_n6992_;
   wire new_n6991_;
   wire new_n6990_1_;
   wire new_n6989_;
   wire new_n6988_;
   wire new_n6987_;
   wire new_n6986_1_;
   wire new_n6985_;
   wire new_n6984_;
   wire new_n6983_;
   wire new_n6982_1_;
   wire new_n6981_;
   wire new_n6980_;
   wire new_n6979_;
   wire new_n6978_;
   wire new_n6977_1_;
   wire new_n6976_;
   wire new_n6975_;
   wire new_n6974_1_;
   wire new_n6973_;
   wire new_n6972_;
   wire new_n6971_;
   wire new_n6970_;
   wire new_n6969_1_;
   wire new_n6968_;
   wire new_n6967_;
   wire new_n6966_;
   wire new_n6965_;
   wire new_n6963_;
   wire new_n6961_;
   wire new_n6960_1_;
   wire new_n6959_;
   wire new_n6957_1_;
   wire new_n6956_;
   wire new_n6955_;
   wire new_n6954_;
   wire new_n6953_;
   wire new_n6952_1_;
   wire new_n6951_;
   wire new_n6950_;
   wire new_n6949_;
   wire new_n6948_;
   wire new_n6947_1_;
   wire new_n6946_;
   wire new_n6945_;
   wire new_n6944_;
   wire new_n6943_1_;
   wire new_n6942_;
   wire new_n6941_;
   wire new_n6940_;
   wire new_n6939_;
   wire new_n6937_;
   wire new_n6936_;
   wire new_n6935_;
   wire new_n6934_1_;
   wire new_n6933_;
   wire new_n6932_;
   wire new_n6920_;
   wire new_n6919_1_;
   wire new_n6918_;
   wire new_n6917_;
   wire new_n6916_;
   wire new_n6915_1_;
   wire new_n6914_;
   wire new_n6913_;
   wire new_n6912_;
   wire new_n6911_;
   wire new_n6910_1_;
   wire new_n6909_;
   wire new_n6907_;
   wire new_n6906_1_;
   wire new_n6905_;
   wire new_n6904_;
   wire new_n6903_;
   wire new_n6902_1_;
   wire new_n6901_;
   wire new_n6900_;
   wire new_n6899_1_;
   wire new_n6898_;
   wire new_n6897_;
   wire new_n6896_;
   wire new_n6895_1_;
   wire new_n6894_;
   wire new_n6893_;
   wire new_n6892_;
   wire new_n6891_;
   wire new_n6890_1_;
   wire new_n6889_;
   wire new_n6888_;
   wire new_n6887_;
   wire new_n6886_1_;
   wire new_n6882_;
   wire new_n6881_1_;
   wire new_n6880_;
   wire new_n6879_;
   wire new_n6878_;
   wire new_n6877_;
   wire new_n6876_1_;
   wire new_n6875_;
   wire new_n6874_;
   wire new_n6873_;
   wire new_n6872_1_;
   wire new_n6871_;
   wire new_n6870_;
   wire new_n6869_;
   wire new_n6868_;
   wire new_n6867_1_;
   wire new_n6866_;
   wire new_n6865_;
   wire new_n6864_;
   wire new_n6863_1_;
   wire new_n6862_;
   wire new_n6861_;
   wire new_n6860_1_;
   wire new_n6859_;
   wire new_n6858_;
   wire new_n6857_;
   wire new_n6856_;
   wire new_n6855_1_;
   wire new_n6854_;
   wire new_n6853_;
   wire new_n6852_;
   wire new_n6851_;
   wire new_n6850_1_;
   wire new_n6849_;
   wire new_n6848_;
   wire new_n6847_;
   wire new_n6846_;
   wire new_n6845_1_;
   wire new_n6844_;
   wire new_n6843_;
   wire new_n6842_;
   wire new_n6841_;
   wire new_n6840_1_;
   wire new_n6839_;
   wire new_n6838_;
   wire new_n6837_;
   wire new_n6836_1_;
   wire new_n6835_;
   wire new_n6834_;
   wire new_n6833_;
   wire new_n6832_;
   wire new_n6831_1_;
   wire new_n6830_;
   wire new_n6829_;
   wire new_n6828_;
   wire new_n6827_;
   wire new_n6826_1_;
   wire new_n6825_;
   wire new_n6823_;
   wire new_n6822_1_;
   wire new_n6821_;
   wire new_n6820_;
   wire new_n6819_;
   wire new_n6815_;
   wire new_n6814_;
   wire new_n6813_1_;
   wire new_n6812_;
   wire new_n6811_;
   wire new_n6810_;
   wire new_n6809_1_;
   wire new_n6808_;
   wire new_n6807_;
   wire new_n6806_1_;
   wire new_n6805_;
   wire new_n6804_;
   wire new_n6803_;
   wire new_n6802_;
   wire new_n6801_1_;
   wire new_n6800_;
   wire new_n6799_;
   wire new_n6798_;
   wire new_n6797_;
   wire new_n6796_1_;
   wire new_n6795_;
   wire new_n6794_;
   wire new_n6793_1_;
   wire new_n6792_;
   wire new_n6791_;
   wire new_n6790_;
   wire new_n6789_;
   wire new_n6788_1_;
   wire new_n6787_;
   wire new_n6786_;
   wire new_n6785_;
   wire new_n6784_;
   wire new_n6783_1_;
   wire new_n6782_;
   wire new_n6781_;
   wire new_n6780_;
   wire new_n6779_1_;
   wire new_n6778_;
   wire new_n6777_;
   wire new_n6776_;
   wire new_n6775_;
   wire new_n6774_1_;
   wire new_n6773_;
   wire new_n6772_;
   wire new_n6771_;
   wire new_n6770_1_;
   wire new_n6769_;
   wire new_n6768_;
   wire new_n6767_;
   wire new_n6766_;
   wire new_n6765_1_;
   wire new_n6764_;
   wire new_n6763_;
   wire new_n6762_;
   wire new_n6761_1_;
   wire new_n6760_;
   wire new_n6759_;
   wire new_n6756_1_;
   wire new_n6755_;
   wire new_n6754_;
   wire new_n6752_1_;
   wire new_n6751_;
   wire new_n6750_;
   wire new_n6749_1_;
   wire new_n6748_;
   wire new_n6747_;
   wire new_n6746_1_;
   wire new_n6745_;
   wire new_n6744_;
   wire new_n6743_;
   wire new_n6742_;
   wire new_n6741_1_;
   wire new_n12336_;
   wire new_n12332_;
   wire new_n12331_;
   wire new_n12330_;
   wire new_n12329_;
   wire new_n12328_;
   wire new_n12327_;
   wire new_n12326_;
   wire new_n12325_;
   wire new_n12324_;
   wire new_n12321_;
   wire new_n12317_;
   wire new_n12316_;
   wire new_n12311_;
   wire new_n12309_;
   wire new_n12308_;
   wire new_n12306_;
   wire new_n12305_;
   wire new_n12304_;
   wire new_n12303_;
   wire new_n12302_;
   wire new_n12301_;
   wire new_n12300_;
   wire new_n12299_;
   wire new_n12298_;
   wire new_n12296_;
   wire new_n12295_;
   wire new_n12294_;
   wire new_n12293_;
   wire new_n12291_;
   wire new_n12290_;
   wire new_n12289_;
   wire new_n12287_;
   wire new_n12286_;
   wire new_n12283_;
   wire new_n12282_;
   wire new_n12281_;
   wire new_n12280_;
   wire new_n12279_;
   wire new_n12278_;
   wire new_n12277_;
   wire new_n12276_;
   wire new_n12275_;
   wire new_n12274_;
   wire new_n12273_;
   wire new_n12272_;
   wire new_n12271_;
   wire new_n12269_;
   wire new_n12266_;
   wire new_n12249_;
   wire new_n12246_;
   wire new_n12245_;
   wire new_n12244_;
   wire new_n12243_;
   wire new_n12242_;
   wire new_n12241_;
   wire new_n12240_;
   wire new_n12239_;
   wire new_n12238_;
   wire new_n12236_;
   wire new_n12235_;
   wire new_n12230_;
   wire new_n12227_;
   wire new_n12218_;
   wire new_n12217_;
   wire new_n12216_;
   wire new_n12215_;
   wire new_n12214_;
   wire new_n12213_;
   wire new_n12212_;
   wire new_n12211_;
   wire new_n12210_;
   wire new_n12209_;
   wire new_n12205_;
   wire new_n12204_;
   wire new_n12202_;
   wire new_n12201_;
   wire new_n12200_;
   wire new_n12199_;
   wire new_n12196_;
   wire new_n12195_;
   wire new_n12190_;
   wire new_n12188_;
   wire new_n12185_;
   wire new_n12184_;
   wire new_n12177_;
   wire new_n12176_;
   wire new_n12175_;
   wire new_n12174_;
   wire new_n12172_;
   wire new_n12170_;
   wire new_n12166_;
   wire new_n12165_;
   wire new_n12164_;
   wire new_n12163_;
   wire new_n12162_;
   wire new_n12155_;
   wire new_n12148_;
   wire new_n12145_;
   wire new_n12141_;
   wire new_n12140_;
   wire new_n12139_;
   wire new_n12138_;
   wire new_n12137_;
   wire new_n12136_;
   wire new_n12135_;
   wire new_n12134_;
   wire new_n12133_;
   wire new_n12131_;
   wire new_n12130_;
   wire new_n12129_;
   wire new_n12128_;
   wire new_n12127_;
   wire new_n12126_;
   wire new_n12125_;
   wire new_n12124_;
   wire new_n12123_;
   wire new_n12122_;
   wire new_n12121_;
   wire new_n12120_;
   wire new_n12119_;
   wire new_n12118_;
   wire new_n12114_;
   wire new_n12113_;
   wire new_n12112_;
   wire new_n12111_;
   wire new_n12110_;
   wire new_n12109_;
   wire new_n12103_;
   wire new_n12097_;
   wire new_n12096_;
   wire new_n12091_;
   wire new_n12090_;
   wire new_n12088_;
   wire new_n12087_;
   wire new_n12079_;
   wire new_n12078_;
   wire new_n12076_;
   wire new_n12075_;
   wire new_n12074_;
   wire new_n12073_;
   wire new_n12072_;
   wire new_n12071_;
   wire new_n12070_;
   wire new_n12069_;
   wire new_n12068_;
   wire new_n12065_;
   wire new_n12061_;
   wire new_n12057_;
   wire new_n12056_;
   wire new_n12053_;
   wire new_n12052_;
   wire new_n12051_;
   wire new_n12050_;
   wire new_n12049_;
   wire new_n12048_;
   wire new_n12047_;
   wire new_n12046_;
   wire new_n12045_;
   wire new_n12044_;
   wire new_n12043_;
   wire new_n12042_;
   wire new_n12041_;
   wire new_n12040_;
   wire new_n12039_;
   wire new_n12038_;
   wire new_n12037_;
   wire new_n12036_;
   wire new_n12035_;
   wire new_n12031_;
   wire new_n12030_;
   wire new_n12020_;
   wire new_n12018_;
   wire new_n12017_;
   wire new_n12008_;
   wire new_n12007_;
   wire new_n12006_;
   wire new_n12005_;
   wire new_n12004_;
   wire new_n12000_;
   wire new_n11999_;
   wire new_n11998_;
   wire new_n11997_;
   wire new_n11996_;
   wire new_n11995_;
   wire new_n11994_;
   wire new_n11993_;
   wire new_n11992_;
   wire new_n11991_;
   wire new_n11990_;
   wire new_n11989_;
   wire new_n11987_;
   wire new_n11982_;
   wire new_n11981_;
   wire new_n11979_;
   wire new_n11978_;
   wire new_n11962_;
   wire new_n11957_;
   wire new_n11953_;
   wire new_n11952_;
   wire new_n11948_;
   wire new_n11941_;
   wire new_n11940_;
   wire new_n11939_;
   wire new_n11938_;
   wire new_n11937_;
   wire new_n11936_;
   wire new_n11935_;
   wire new_n11934_;
   wire new_n11933_;
   wire new_n11931_;
   wire new_n11930_;
   wire new_n11928_;
   wire new_n11927_;
   wire new_n11924_;
   wire new_n11922_;
   wire new_n11912_;
   wire new_n11911_;
   wire new_n11910_;
   wire new_n11909_;
   wire new_n11908_;
   wire new_n11907_;
   wire new_n11906_;
   wire new_n11905_;
   wire new_n11904_;
   wire new_n11901_;
   wire new_n11898_;
   wire new_n11895_;
   wire new_n11893_;
   wire new_n11892_;
   wire new_n11884_;
   wire new_n11883_;
   wire new_n11881_;
   wire new_n11868_;
   wire new_n11867_;
   wire new_n11856_;
   wire new_n11855_;
   wire new_n11852_;
   wire new_n11851_;
   wire new_n11847_;
   wire new_n11846_;
   wire new_n11845_;
   wire new_n11844_;
   wire new_n11843_;
   wire new_n11842_;
   wire new_n11841_;
   wire new_n11840_;
   wire new_n11839_;
   wire new_n11832_;
   wire new_n11831_;
   wire new_n11829_;
   wire new_n11823_;
   wire new_n11820_;
   wire new_n11816_;
   wire new_n11815_;
   wire new_n11813_;
   wire new_n11812_;
   wire new_n11805_;
   wire new_n11803_;
   wire new_n11802_;
   wire new_n11787_;
   wire new_n11785_;
   wire new_n11784_;
   wire new_n11780_;
   wire new_n11776_;
   wire new_n11775_;
   wire new_n11772_;
   wire new_n11764_;
   wire new_n11763_;
   wire new_n11761_;
   wire new_n11760_;
   wire new_n11759_;
   wire new_n11758_;
   wire new_n11757_;
   wire new_n11755_;
   wire new_n11749_;
   wire new_n11744_;
   wire new_n11743_;
   wire new_n11742_;
   wire new_n11741_;
   wire new_n11739_;
   wire new_n11738_;
   wire new_n11736_;
   wire new_n11732_;
   wire new_n11731_;
   wire new_n11730_;
   wire new_n11729_;
   wire new_n11728_;
   wire new_n11727_;
   wire new_n11726_;
   wire new_n11725_;
   wire new_n11724_;
   wire new_n11723_;
   wire new_n11722_;
   wire new_n11721_;
   wire new_n11720_;
   wire new_n11716_;
   wire new_n11715_;
   wire new_n11709_;
   wire new_n11708_;
   wire new_n11705_;
   wire new_n11700_;
   wire new_n11699_;
   wire new_n11698_;
   wire new_n11697_;
   wire new_n11696_;
   wire new_n11695_;
   wire new_n11694_;
   wire new_n11693_;
   wire new_n11692_;
   wire new_n11686_;
   wire new_n11683_;
   wire new_n11680_;
   wire new_n11679_;
   wire new_n11678_;
   wire new_n11676_;
   wire new_n11675_;
   wire new_n11671_;
   wire new_n11663_;
   wire new_n11662_;
   wire new_n11657_;
   wire new_n11656_;
   wire new_n11653_;
   wire new_n11651_;
   wire new_n11646_;
   wire new_n11640_;
   wire new_n11639_;
   wire new_n11638_;
   wire new_n11637_;
   wire new_n11636_;
   wire new_n11635_;
   wire new_n11634_;
   wire new_n11633_;
   wire new_n11632_;
   wire new_n11631_;
   wire new_n11630_;
   wire new_n11629_;
   wire new_n11628_;
   wire new_n11627_;
   wire new_n11625_;
   wire new_n11624_;
   wire new_n11613_;
   wire new_n11612_;
   wire new_n11611_;
   wire new_n11610_;
   wire new_n11609_;
   wire new_n11608_;
   wire new_n11607_;
   wire new_n11606_;
   wire new_n11605_;
   wire new_n11604_;
   wire new_n11601_;
   wire new_n11600_;
   wire new_n11599_;
   wire new_n11598_;
   wire new_n11593_;
   wire new_n11592_;
   wire new_n11590_;
   wire new_n11589_;
   wire new_n11584_;
   wire new_n11583_;
   wire new_n11582_;
   wire new_n11581_;
   wire new_n11578_;
   wire new_n11576_;
   wire new_n11575_;
   wire new_n11574_;
   wire new_n11573_;
   wire new_n11568_;
   wire new_n11567_;
   wire new_n11564_;
   wire new_n11563_;
   wire new_n11562_;
   wire new_n11561_;
   wire new_n11560_;
   wire new_n11559_;
   wire new_n11558_;
   wire new_n11557_;
   wire new_n11556_;
   wire new_n11555_;
   wire new_n11554_;
   wire new_n11553_;
   wire new_n11552_;
   wire new_n11551_;
   wire new_n11550_;
   wire new_n11535_;
   wire new_n11534_;
   wire new_n11527_;
   wire new_n11525_;
   wire new_n11524_;
   wire new_n11513_;
   wire new_n11512_;
   wire new_n11509_;
   wire new_n11508_;
   wire new_n11507_;
   wire new_n11506_;
   wire new_n11505_;
   wire new_n11504_;
   wire new_n11503_;
   wire new_n11502_;
   wire new_n11501_;
   wire new_n11499_;
   wire new_n11498_;
   wire new_n11494_;
   wire new_n11493_;
   wire new_n11492_;
   wire new_n11489_;
   wire new_n11488_;
   wire new_n11485_;
   wire new_n11484_;
   wire new_n11481_;
   wire new_n11475_;
   wire new_n11470_;
   wire new_n11469_;
   wire new_n11468_;
   wire new_n11467_;
   wire new_n11466_;
   wire new_n11465_;
   wire new_n11464_;
   wire new_n11463_;
   wire new_n11462_;
   wire new_n11461_;
   wire new_n11459_;
   wire new_n11458_;
   wire new_n11456_;
   wire new_n11455_;
   wire new_n11449_;
   wire new_n11448_;
   wire new_n11436_;
   wire new_n11435_;
   wire new_n11434_;
   wire new_n11433_;
   wire new_n11432_;
   wire new_n11431_;
   wire new_n11430_;
   wire new_n11429_;
   wire new_n11428_;
   wire new_n11422_;
   wire new_n11421_;
   wire new_n11419_;
   wire new_n11418_;
   wire new_n11417_;
   wire new_n11416_;
   wire new_n11409_;
   wire new_n11408_;
   wire new_n11406_;
   wire new_n11405_;
   wire new_n11404_;
   wire new_n11402_;
   wire new_n11395_;
   wire new_n11394_;
   wire new_n11389_;
   wire new_n11388_;
   wire new_n11382_;
   wire new_n11381_;
   wire new_n11377_;
   wire new_n11374_;
   wire new_n11367_;
   wire new_n11364_;
   wire new_n11363_;
   wire new_n11360_;
   wire new_n11359_;
   wire new_n11358_;
   wire new_n11357_;
   wire new_n11356_;
   wire new_n11355_;
   wire new_n11354_;
   wire new_n11353_;
   wire new_n11350_;
   wire new_n11349_;
   wire new_n11345_;
   wire new_n11344_;
   wire new_n11337_;
   wire new_n11336_;
   wire new_n11334_;
   wire new_n11333_;
   wire new_n11332_;
   wire new_n11330_;
   wire new_n11329_;
   wire new_n11328_;
   wire new_n11327_;
   wire new_n11326_;
   wire new_n11325_;
   wire new_n11324_;
   wire new_n11323_;
   wire new_n11322_;
   wire new_n11317_;
   wire new_n11316_;
   wire new_n11315_;
   wire new_n11314_;
   wire new_n11313_;
   wire new_n11312_;
   wire new_n11311_;
   wire new_n11310_;
   wire new_n11309_;
   wire new_n11308_;
   wire new_n11301_;
   wire new_n11298_;
   wire new_n11297_;
   wire new_n11296_;
   wire new_n11295_;
   wire new_n11294_;
   wire new_n11293_;
   wire new_n11292_;
   wire new_n11291_;
   wire new_n11290_;
   wire new_n11289_;
   wire new_n11288_;
   wire new_n11287_;
   wire new_n11286_;
   wire new_n11285_;
   wire new_n11282_;
   wire new_n11280_;
   wire new_n11279_;
   wire new_n11271_;
   wire new_n11270_;
   wire new_n11267_;
   wire new_n11266_;
   wire new_n11265_;
   wire new_n11264_;
   wire new_n11263_;
   wire new_n11262_;
   wire new_n11261_;
   wire new_n11260_;
   wire new_n11259_;
   wire new_n11257_;
   wire new_n11256_;
   wire new_n11255_;
   wire new_n11254_;
   wire new_n11253_;
   wire new_n11252_;
   wire new_n11251_;
   wire new_n11250_;
   wire new_n11249_;
   wire new_n11248_;
   wire new_n11247_;
   wire new_n11246_;
   wire new_n11244_;
   wire new_n11243_;
   wire new_n11242_;
   wire new_n11233_;
   wire new_n11232_;
   wire new_n11227_;
   wire new_n11225_;
   wire new_n11221_;
   wire new_n11220_;
   wire new_n11214_;
   wire new_n11213_;
   wire new_n11210_;
   wire new_n11208_;
   wire new_n11207_;
   wire new_n11206_;
   wire new_n11205_;
   wire new_n11202_;
   wire new_n11201_;
   wire new_n11199_;
   wire new_n11198_;
   wire new_n11197_;
   wire new_n11195_;
   wire new_n11194_;
   wire new_n11193_;
   wire new_n11192_;
   wire new_n11191_;
   wire new_n11190_;
   wire new_n11189_;
   wire new_n11188_;
   wire new_n11187_;
   wire new_n11186_;
   wire new_n11185_;
   wire new_n11184_;
   wire new_n11183_;
   wire new_n11182_;
   wire new_n11176_;
   wire new_n11175_;
   wire new_n11169_;
   wire new_n11168_;
   wire new_n11167_;
   wire new_n11166_;
   wire new_n11163_;
   wire new_n11160_;
   wire new_n11155_;
   wire new_n11154_;
   wire new_n11148_;
   wire new_n11147_;
   wire new_n11146_;
   wire new_n11145_;
   wire new_n11141_;
   wire new_n11140_;
   wire new_n11134_;
   wire new_n11130_;
   wire new_n11129_;
   wire new_n11123_;
   wire new_n11122_;
   wire new_n11121_;
   wire new_n11118_;
   wire new_n11117_;
   wire new_n11113_;
   wire new_n11112_;
   wire new_n11111_;
   wire new_n11110_;
   wire new_n11109_;
   wire new_n11108_;
   wire new_n11107_;
   wire new_n11106_;
   wire new_n11105_;
   wire new_n11100_;
   wire new_n11090_;
   wire new_n11087_;
   wire new_n11086_;
   wire new_n11085_;
   wire new_n11084_;
   wire new_n11077_;
   wire new_n11076_;
   wire new_n11074_;
   wire new_n11073_;
   wire new_n11067_;
   wire new_n11064_;
   wire new_n11063_;
   wire new_n11062_;
   wire new_n11061_;
   wire new_n11060_;
   wire new_n11059_;
   wire new_n11058_;
   wire new_n11057_;
   wire new_n11056_;
   wire new_n11052_;
   wire new_n11047_;
   wire new_n11046_;
   wire new_n11045_;
   wire new_n11041_;
   wire new_n11040_;
   wire new_n11039_;
   wire new_n11038_;
   wire new_n11037_;
   wire new_n11036_;
   wire new_n11035_;
   wire new_n11034_;
   wire new_n11027_;
   wire new_n11019_;
   wire new_n11018_;
   wire new_n11017_;
   wire new_n11015_;
   wire new_n11006_;
   wire new_n11005_;
   wire new_n11004_;
   wire new_n11003_;
   wire new_n11002_;
   wire new_n11001_;
   wire new_n11000_;
   wire new_n10999_;
   wire new_n10998_;
   wire new_n10997_;
   wire new_n10994_;
   wire new_n10993_;
   wire new_n10986_;
   wire new_n10985_;
   wire new_n10982_;
   wire new_n10981_;
   wire new_n10979_;
   wire new_n10978_;
   wire new_n10977_;
   wire new_n10976_;
   wire new_n10975_;
   wire new_n10974_;
   wire new_n10973_;
   wire new_n10972_;
   wire new_n10971_;
   wire new_n10969_;
   wire new_n10968_;
   wire new_n10963_;
   wire new_n10962_;
   wire new_n10955_;
   wire new_n10954_;
   wire new_n10952_;
   wire new_n10951_;
   wire new_n10950_;
   wire new_n10949_;
   wire new_n10948_;
   wire new_n10947_;
   wire new_n10946_;
   wire new_n10945_;
   wire new_n10944_;
   wire new_n10940_;
   wire new_n10939_;
   wire new_n10933_;
   wire new_n10932_;
   wire new_n10930_;
   wire new_n10929_;
   wire new_n10926_;
   wire new_n10925_;
   wire new_n10918_;
   wire new_n10917_;
   wire new_n10914_;
   wire new_n10913_;
   wire new_n10912_;
   wire new_n10911_;
   wire new_n10910_;
   wire new_n10909_;
   wire new_n10908_;
   wire new_n10907_;
   wire new_n10906_;
   wire new_n10903_;
   wire new_n10902_;
   wire new_n10896_;
   wire new_n10895_;
   wire new_n10893_;
   wire new_n10892_;
   wire new_n10890_;
   wire new_n10880_;
   wire new_n10879_;
   wire new_n10875_;
   wire new_n10874_;
   wire new_n10871_;
   wire new_n10869_;
   wire new_n10868_;
   wire new_n10867_;
   wire new_n10866_;
   wire new_n10865_;
   wire new_n10864_;
   wire new_n10863_;
   wire new_n10862_;
   wire new_n10861_;
   wire new_n10860_;
   wire new_n10857_;
   wire new_n10856_;
   wire new_n10855_;
   wire new_n10854_;
   wire new_n10853_;
   wire new_n10852_;
   wire new_n10851_;
   wire new_n10850_;
   wire new_n10849_;
   wire new_n10839_;
   wire new_n10838_;
   wire new_n10837_;
   wire new_n10836_;
   wire new_n10835_;
   wire new_n10834_;
   wire new_n10833_;
   wire new_n10832_;
   wire new_n10831_;
   wire new_n10830_;
   wire new_n10829_;
   wire new_n10828_;
   wire new_n10827_;
   wire new_n10826_;
   wire new_n10825_;
   wire new_n10824_;
   wire new_n10823_;
   wire new_n10822_;
   wire new_n10821_;
   wire new_n10820_;
   wire new_n10819_;
   wire new_n10818_;
   wire new_n10817_;
   wire new_n10816_;
   wire new_n10815_;
   wire new_n10811_;
   wire new_n10810_;
   wire new_n10805_;
   wire new_n10804_;
   wire new_n10803_;
   wire new_n10802_;
   wire new_n10801_;
   wire new_n10800_;
   wire new_n10799_;
   wire new_n10798_;
   wire new_n10797_;
   wire new_n10796_;
   wire new_n10795_;
   wire new_n10794_;
   wire new_n10793_;
   wire new_n10792_;
   wire new_n10785_;
   wire new_n10784_;
   wire new_n10783_;
   wire new_n10782_;
   wire new_n10781_;
   wire new_n10780_;
   wire new_n10779_;
   wire new_n10778_;
   wire new_n10777_;
   wire new_n10776_;
   wire new_n10775_;
   wire new_n10774_;
   wire new_n10767_;
   wire new_n10766_;
   wire new_n10765_;
   wire new_n10764_;
   wire new_n10761_;
   wire new_n10756_;
   wire new_n10755_;
   wire new_n10754_;
   wire new_n10753_;
   wire new_n10752_;
   wire new_n10751_;
   wire new_n10749_;
   wire new_n10748_;
   wire new_n10746_;
   wire new_n10745_;
   wire new_n10744_;
   wire new_n10743_;
   wire new_n10742_;
   wire new_n10741_;
   wire new_n10740_;
   wire new_n10739_;
   wire new_n10738_;
   wire new_n10737_;
   wire new_n10736_;
   wire new_n10735_;
   wire new_n10734_;
   wire new_n10733_;
   wire new_n10732_;
   wire new_n10730_;
   wire new_n10729_;
   wire new_n10726_;
   wire new_n10725_;
   wire new_n10721_;
   wire new_n10720_;
   wire new_n10712_;
   wire new_n10711_;
   wire new_n10707_;
   wire new_n10706_;
   wire new_n10704_;
   wire new_n10703_;
   wire new_n10702_;
   wire new_n10701_;
   wire new_n10692_;
   wire new_n10691_;
   wire new_n10690_;
   wire new_n10680_;
   wire new_n10679_;
   wire new_n10677_;
   wire new_n10673_;
   wire new_n10672_;
   wire new_n10666_;
   wire new_n10665_;
   wire new_n10660_;
   wire new_n10659_;
   wire new_n10658_;
   wire new_n10657_;
   wire new_n10656_;
   wire new_n10655_;
   wire new_n10654_;
   wire new_n10653_;
   wire new_n10652_;
   wire new_n10651_;
   wire new_n10650_;
   wire new_n10649_;
   wire new_n10648_;
   wire new_n10647_;
   wire new_n10642_;
   wire new_n10641_;
   wire new_n10640_;
   wire new_n10637_;
   wire new_n10636_;
   wire new_n10631_;
   wire new_n10628_;
   wire new_n10627_;
   wire new_n10626_;
   wire new_n10625_;
   wire new_n10624_;
   wire new_n10623_;
   wire new_n10622_;
   wire new_n10621_;
   wire new_n10620_;
   wire new_n10619_;
   wire new_n10618_;
   wire new_n10617_;
   wire new_n10616_;
   wire new_n10615_;
   wire new_n10608_;
   wire new_n10607_;
   wire new_n10606_;
   wire new_n10605_;
   wire new_n10600_;
   wire new_n10599_;
   wire new_n10598_;
   wire new_n10597_;
   wire new_n10595_;
   wire new_n10594_;
   wire new_n10593_;
   wire new_n10592_;
   wire new_n10591_;
   wire new_n10590_;
   wire new_n10589_;
   wire new_n10588_;
   wire new_n10587_;
   wire new_n10586_;
   wire new_n10585_;
   wire new_n10584_;
   wire new_n10583_;
   wire new_n10582_;
   wire new_n10579_;
   wire new_n10576_;
   wire new_n10575_;
   wire new_n10573_;
   wire new_n10572_;
   wire new_n10567_;
   wire new_n10566_;
   wire new_n10564_;
   wire new_n10559_;
   wire new_n10558_;
   wire new_n10557_;
   wire new_n10556_;
   wire new_n10555_;
   wire new_n10552_;
   wire new_n10551_;
   wire new_n10550_;
   wire new_n10549_;
   wire new_n10548_;
   wire new_n10547_;
   wire new_n10546_;
   wire new_n10545_;
   wire new_n10544_;
   wire new_n10543_;
   wire new_n10542_;
   wire new_n10541_;
   wire new_n10540_;
   wire new_n10539_;
   wire new_n10536_;
   wire new_n10535_;
   wire new_n10530_;
   wire new_n10529_;
   wire new_n10528_;
   wire new_n10527_;
   wire new_n10526_;
   wire new_n10525_;
   wire new_n10524_;
   wire new_n10522_;
   wire new_n10521_;
   wire new_n10517_;
   wire new_n10516_;
   wire new_n10515_;
   wire new_n10514_;
   wire new_n10506_;
   wire new_n10505_;
   wire new_n10499_;
   wire new_n10498_;
   wire new_n10497_;
   wire new_n10496_;
   wire new_n10495_;
   wire new_n10494_;
   wire new_n10493_;
   wire new_n10492_;
   wire new_n10491_;
   wire new_n10490_;
   wire new_n10489_;
   wire new_n10488_;
   wire new_n10487_;
   wire new_n10486_;
   wire new_n10479_;
   wire new_n10478_;
   wire new_n10476_;
   wire new_n10475_;
   wire new_n10473_;
   wire new_n10472_;
   wire new_n10469_;
   wire new_n10468_;
   wire new_n10464_;
   wire new_n10463_;
   wire new_n10460_;
   wire new_n10459_;
   wire new_n10458_;
   wire new_n10457_;
   wire new_n10456_;
   wire new_n10455_;
   wire new_n10454_;
   wire new_n10453_;
   wire new_n10452_;
   wire new_n10448_;
   wire new_n10447_;
   wire new_n10444_;
   wire new_n10443_;
   wire new_n10442_;
   wire new_n10441_;
   wire new_n10440_;
   wire new_n10439_;
   wire new_n10438_;
   wire new_n10437_;
   wire new_n10436_;
   wire new_n10428_;
   wire new_n10427_;
   wire new_n10425_;
   wire new_n10424_;
   wire new_n10422_;
   wire new_n10421_;
   wire new_n10419_;
   wire new_n10418_;
   wire new_n10417_;
   wire new_n10414_;
   wire new_n10413_;
   wire new_n10395_;
   wire new_n10394_;
   wire new_n10390_;
   wire new_n10389_;
   wire new_n10380_;
   wire new_n10379_;
   wire new_n10377_;
   wire new_n10376_;
   wire new_n10371_;
   wire new_n10368_;
   wire new_n10367_;
   wire new_n10364_;
   wire new_n10359_;
   wire new_n10354_;
   wire new_n10353_;
   wire new_n10352_;
   wire new_n10351_;
   wire new_n10350_;
   wire new_n10349_;
   wire new_n10348_;
   wire new_n10347_;
   wire new_n10346_;
   wire new_n10340_;
   wire new_n10339_;
   wire new_n10337_;
   wire new_n10336_;
   wire new_n10335_;
   wire new_n10325_;
   wire new_n10322_;
   wire new_n10314_;
   wire new_n10305_;
   wire new_n10303_;
   wire new_n10302_;
   wire new_n10301_;
   wire new_n10300_;
   wire new_n10299_;
   wire new_n10298_;
   wire new_n10297_;
   wire new_n10296_;
   wire new_n10295_;
   wire new_n10294_;
   wire new_n10293_;
   wire new_n10292_;
   wire new_n10291_;
   wire new_n10290_;
   wire new_n10284_;
   wire new_n10283_;
   wire new_n10281_;
   wire new_n10280_;
   wire new_n10279_;
   wire new_n10278_;
   wire new_n10277_;
   wire new_n10276_;
   wire new_n10275_;
   wire new_n10274_;
   wire new_n10273_;
   wire new_n10266_;
   wire new_n10265_;
   wire new_n10263_;
   wire new_n10262_;
   wire new_n10253_;
   wire new_n10252_;
   wire new_n10250_;
   wire new_n10249_;
   wire new_n10248_;
   wire new_n10247_;
   wire new_n10246_;
   wire new_n10245_;
   wire new_n10244_;
   wire new_n10242_;
   wire new_n10241_;
   wire new_n10240_;
   wire new_n10239_;
   wire new_n10238_;
   wire new_n10237_;
   wire new_n10234_;
   wire new_n10233_;
   wire new_n10232_;
   wire new_n10231_;
   wire new_n10230_;
   wire new_n10229_;
   wire new_n10228_;
   wire new_n10227_;
   wire new_n10226_;
   wire new_n10225_;
   wire new_n10222_;
   wire new_n10221_;
   wire new_n10216_;
   wire new_n10215_;
   wire new_n10198_;
   wire new_n10197_;
   wire new_n10193_;
   wire new_n10192_;
   wire new_n10189_;
   wire new_n10188_;
   wire new_n10185_;
   wire new_n10184_;
   wire new_n10183_;
   wire new_n10182_;
   wire new_n10181_;
   wire new_n10180_;
   wire new_n10179_;
   wire new_n10178_;
   wire new_n10177_;
   wire new_n10176_;
   wire new_n10175_;
   wire new_n10174_;
   wire new_n10173_;
   wire new_n10172_;
   wire new_n10163_;
   wire new_n10162_;
   wire new_n10159_;
   wire new_n10158_1_;
   wire new_n10157_;
   wire new_n10151_;
   wire new_n10150_1_;
   wire new_n10148_;
   wire new_n10147_;
   wire new_n10144_;
   wire new_n10143_;
   wire new_n10136_;
   wire new_n10135_;
   wire new_n10133_;
   wire new_n10132_1_;
   wire new_n10131_;
   wire new_n10130_;
   wire new_n10129_;
   wire new_n10126_;
   wire new_n10125_;
   wire new_n10121_;
   wire new_n10115_;
   wire new_n10114_;
   wire new_n10112_1_;
   wire new_n10111_;
   wire new_n10110_;
   wire new_n10106_;
   wire new_n10105_;
   wire new_n10104_;
   wire new_n10103_1_;
   wire new_n10102_;
   wire new_n10101_;
   wire new_n10100_;
   wire new_n10099_1_;
   wire new_n10098_;
   wire new_n10097_;
   wire new_n10095_;
   wire new_n10094_1_;
   wire new_n10093_;
   wire new_n10092_;
   wire new_n10091_;
   wire new_n10090_;
   wire new_n10089_1_;
   wire new_n10086_;
   wire new_n10085_;
   wire new_n10084_1_;
   wire new_n10076_;
   wire new_n10075_;
   wire new_n10068_;
   wire new_n10067_;
   wire new_n10064_;
   wire new_n10063_;
   wire new_n10058_;
   wire new_n10056_1_;
   wire new_n10055_;
   wire new_n10054_;
   wire new_n10053_;
   wire new_n10052_1_;
   wire new_n10051_;
   wire new_n10049_;
   wire new_n10047_1_;
   wire new_n10046_;
   wire new_n10045_;
   wire new_n10044_;
   wire new_n10043_;
   wire new_n10042_1_;
   wire new_n10041_;
   wire new_n10040_;
   wire new_n10039_;
   wire new_n10038_;
   wire new_n10035_;
   wire new_n10034_;
   wire new_n10031_;
   wire new_n10030_;
   wire new_n10028_1_;
   wire new_n10027_;
   wire new_n10025_;
   wire new_n10021_;
   wire new_n10010_1_;
   wire new_n10009_;
   wire new_n10008_;
   wire new_n10006_1_;
   wire new_n10005_;
   wire net_7807;
   wire net_7802;
   wire net_7799;
   wire net_7792;
   wire net_7790;
   wire net_7780;
   wire net_7779;
   wire net_7778;
   wire net_7777;
   wire net_7776;
   wire net_7775;
   wire net_7774;
   wire net_7773;
   wire net_7772;
   wire net_7771;
   wire net_7770;
   wire net_7769;
   wire net_7767;
   wire net_7766;
   wire net_7764;
   wire net_7762;
   wire net_7760;
   wire net_7758;
   wire net_7756;
   wire net_7754;
   wire net_7752;
   wire net_7750;
   wire net_7744;
   wire net_7743;
   wire net_7742;
   wire net_7741;
   wire net_7740;
   wire net_7739;
   wire net_7738;
   wire net_7737;
   wire net_7715;
   wire net_7714;
   wire net_7713;
   wire net_7712;
   wire net_7711;
   wire net_7710;
   wire net_7709;
   wire net_7708;
   wire net_7691;
   wire net_7680;
   wire net_7679;
   wire net_7678;
   wire net_7677;
   wire net_7676;
   wire net_7675;
   wire net_7674;
   wire net_7673;
   wire net_7672;
   wire net_7671;
   wire net_7670;
   wire net_7669;
   wire net_7668;
   wire net_7647;
   wire net_7646;
   wire net_7645;
   wire net_7644;
   wire net_7643;
   wire net_7642;
   wire net_7641;
   wire net_7640;
   wire net_7639;
   wire net_7638;
   wire net_7637;
   wire net_7636;
   wire net_7615;
   wire net_7614;
   wire net_7613;
   wire net_7612;
   wire net_7611;
   wire net_7610;
   wire net_7609;
   wire net_7608;
   wire net_7607;
   wire net_7606;
   wire net_7605;
   wire net_7604;
   wire net_7551;
   wire net_7550;
   wire net_7549;
   wire net_7548;
   wire net_7547;
   wire net_7546;
   wire net_7545;
   wire net_7544;
   wire net_7543;
   wire net_7542;
   wire net_7541;
   wire net_7540;
   wire net_7539;
   wire net_7538;
   wire net_7537;
   wire net_7536;
   wire net_7529;
   wire net_7528;
   wire net_7527;
   wire net_7526;
   wire net_7525;
   wire net_7524;
   wire net_7523;
   wire net_7522;
   wire net_7521;
   wire net_7520;
   wire net_7519;
   wire net_7518;
   wire net_7517;
   wire net_7496;
   wire net_7495;
   wire net_7494;
   wire net_7493;
   wire net_7492;
   wire net_7491;
   wire net_7490;
   wire net_7489;
   wire net_7488;
   wire net_7487;
   wire net_7486;
   wire net_7485;
   wire net_7464;
   wire net_7463;
   wire net_7462;
   wire net_7461;
   wire net_7460;
   wire net_7459;
   wire net_7458;
   wire net_7457;
   wire net_7456;
   wire net_7455;
   wire net_7454;
   wire net_7453;
   wire net_7400;
   wire net_7399;
   wire net_7398;
   wire net_7397;
   wire net_7396;
   wire net_7395;
   wire net_7394;
   wire net_7393;
   wire net_7392;
   wire net_7391;
   wire net_7390;
   wire net_7389;
   wire net_7388;
   wire net_7387;
   wire net_7386;
   wire net_7385;
   wire net_7378;
   wire net_7377;
   wire net_7376;
   wire net_7375;
   wire net_7374;
   wire net_7373;
   wire net_7372;
   wire net_7371;
   wire net_7370;
   wire net_7369;
   wire net_7368;
   wire net_7367;
   wire net_7366;
   wire net_7345;
   wire net_7344;
   wire net_7343;
   wire net_7342;
   wire net_7341;
   wire net_7340;
   wire net_7339;
   wire net_7338;
   wire net_7337;
   wire net_7336;
   wire net_7335;
   wire net_7334;
   wire net_7313;
   wire net_7312;
   wire net_7311;
   wire net_7310;
   wire net_7309;
   wire net_7308;
   wire net_7307;
   wire net_7306;
   wire net_7305;
   wire net_7304;
   wire net_7303;
   wire net_7302;
   wire net_7249;
   wire net_7248;
   wire net_7247;
   wire net_7246;
   wire net_7245;
   wire net_7244;
   wire net_7243;
   wire net_7242;
   wire net_7241;
   wire net_7240;
   wire net_7239;
   wire net_7238;
   wire net_7237;
   wire net_7236;
   wire net_7235;
   wire net_7234;
   wire net_7231;
   wire net_7226;
   wire net_7225;
   wire net_7224;
   wire net_7223;
   wire net_7222;
   wire net_7221;
   wire net_7220;
   wire net_7219;
   wire net_7218;
   wire net_7217;
   wire net_7216;
   wire net_7215;
   wire net_7214;
   wire net_7213;
   wire net_7212;
   wire net_7211;
   wire net_7210;
   wire net_7209;
   wire net_7208;
   wire net_7207;
   wire net_7206;
   wire net_7205;
   wire net_7204;
   wire net_7203;
   wire net_7202;
   wire net_7201;
   wire net_7200;
   wire net_7199;
   wire net_7198;
   wire net_7197;
   wire net_7196;
   wire net_7195;
   wire net_7194;
   wire net_7193;
   wire net_7192;
   wire net_7191;
   wire net_7190;
   wire net_7189;
   wire net_7188;
   wire net_7187;
   wire net_7186;
   wire net_7185;
   wire net_7184;
   wire net_7183;
   wire net_7182;
   wire net_7181;
   wire net_7180;
   wire net_7179;
   wire net_7178;
   wire net_7177;
   wire net_7176;
   wire net_7175;
   wire net_7174;
   wire net_7173;
   wire net_7172;
   wire net_7171;
   wire net_7170;
   wire net_7169;
   wire net_7168;
   wire net_7167;
   wire net_7166;
   wire net_7165;
   wire net_7164;
   wire net_7163;
   wire net_7162;
   wire net_7161;
   wire net_7160;
   wire net_7159;
   wire net_7158;
   wire net_7157;
   wire net_7156;
   wire net_7155;
   wire net_7154;
   wire net_7153;
   wire net_7152;
   wire net_7151;
   wire net_7150;
   wire net_7149;
   wire net_7148;
   wire net_7147;
   wire net_7146;
   wire net_7145;
   wire net_7144;
   wire net_7143;
   wire net_7142;
   wire net_7141;
   wire net_7140;
   wire net_7139;
   wire net_7138;
   wire net_7137;
   wire net_7136;
   wire net_7135;
   wire net_7134;
   wire net_7133;
   wire net_7132;
   wire net_7131;
   wire net_7130;
   wire net_7129;
   wire net_7128;
   wire net_7127;
   wire net_7126;
   wire net_7125;
   wire net_7124;
   wire net_7123;
   wire net_7122;
   wire net_7121;
   wire net_7120;
   wire net_7119;
   wire net_7118;
   wire net_7117;
   wire net_7116;
   wire net_7115;
   wire net_7114;
   wire net_7113;
   wire net_7112;
   wire net_7111;
   wire net_7110;
   wire net_7109;
   wire net_7108;
   wire net_7107;
   wire net_7106;
   wire net_7105;
   wire net_7104;
   wire net_7103;
   wire net_7102;
   wire net_7101;
   wire net_7100;
   wire net_7099;
   wire net_7096;
   wire net_7091;
   wire net_7090;
   wire net_7089;
   wire net_7088;
   wire net_7087;
   wire net_7086;
   wire net_7085;
   wire net_7084;
   wire net_7083;
   wire net_7082;
   wire net_7081;
   wire net_7080;
   wire net_7079;
   wire net_7078;
   wire net_7077;
   wire net_7076;
   wire net_7075;
   wire net_7074;
   wire net_7073;
   wire net_7072;
   wire net_7071;
   wire net_7070;
   wire net_7069;
   wire net_7068;
   wire net_7067;
   wire net_7066;
   wire net_7065;
   wire net_7064;
   wire net_7063;
   wire net_7062;
   wire net_7061;
   wire net_7060;
   wire net_7059;
   wire net_7058;
   wire net_7057;
   wire net_7056;
   wire net_7055;
   wire net_7054;
   wire net_7053;
   wire net_7052;
   wire net_7051;
   wire net_7050;
   wire net_7049;
   wire net_7048;
   wire net_7047;
   wire net_7046;
   wire net_7045;
   wire net_7044;
   wire net_7043;
   wire net_7042;
   wire net_7041;
   wire net_7040;
   wire net_7039;
   wire net_7038;
   wire net_7037;
   wire net_7036;
   wire net_7035;
   wire net_7034;
   wire net_7033;
   wire net_7032;
   wire net_7031;
   wire net_7030;
   wire net_7029;
   wire net_7028;
   wire net_7027;
   wire net_7026;
   wire net_7025;
   wire net_7024;
   wire net_7023;
   wire net_7022;
   wire net_7021;
   wire net_7020;
   wire net_7019;
   wire net_7018;
   wire net_7017;
   wire net_7016;
   wire net_7015;
   wire net_7014;
   wire net_7013;
   wire net_7012;
   wire net_7011;
   wire net_7010;
   wire net_7009;
   wire net_7008;
   wire net_7007;
   wire net_7006;
   wire net_7005;
   wire net_7004;
   wire net_7003;
   wire net_7002;
   wire net_7001;
   wire net_7000;
   wire net_6999;
   wire net_6998;
   wire net_6997;
   wire net_6996;
   wire net_6995;
   wire net_6994;
   wire net_6993;
   wire net_6992;
   wire net_6991;
   wire net_6990;
   wire net_6989;
   wire net_6988;
   wire net_6987;
   wire net_6986;
   wire net_6985;
   wire net_6984;
   wire net_6983;
   wire net_6982;
   wire net_6981;
   wire net_6980;
   wire net_6979;
   wire net_6978;
   wire net_6977;
   wire net_6976;
   wire net_6975;
   wire net_6974;
   wire net_6973;
   wire net_6972;
   wire net_6971;
   wire net_6970;
   wire net_6969;
   wire net_6968;
   wire net_6967;
   wire net_6966;
   wire net_6965;
   wire net_6964;
   wire net_6961;
   wire net_6956;
   wire net_6955;
   wire net_6954;
   wire net_6953;
   wire net_6952;
   wire net_6951;
   wire net_6950;
   wire net_6949;
   wire net_6948;
   wire net_6947;
   wire net_6946;
   wire net_6945;
   wire net_6944;
   wire net_6943;
   wire net_6942;
   wire net_6941;
   wire net_6940;
   wire net_6939;
   wire net_6938;
   wire net_6937;
   wire net_6936;
   wire net_6935;
   wire net_6934;
   wire net_6933;
   wire net_6932;
   wire net_6931;
   wire net_6930;
   wire net_6929;
   wire net_6928;
   wire net_6927;
   wire net_6926;
   wire net_6925;
   wire net_6924;
   wire net_6923;
   wire net_6922;
   wire net_6921;
   wire net_6920;
   wire net_6919;
   wire net_6918;
   wire net_6917;
   wire net_6916;
   wire net_6915;
   wire net_6914;
   wire net_6913;
   wire net_6912;
   wire net_6911;
   wire net_6910;
   wire net_6909;
   wire net_6908;
   wire net_6907;
   wire net_6906;
   wire net_6905;
   wire net_6904;
   wire net_6903;
   wire net_6902;
   wire net_6901;
   wire net_6900;
   wire net_6899;
   wire net_6898;
   wire net_6897;
   wire net_6896;
   wire net_6895;
   wire net_6894;
   wire net_6893;
   wire net_6892;
   wire net_6891;
   wire net_6890;
   wire net_6889;
   wire net_6888;
   wire net_6887;
   wire net_6886;
   wire net_6885;
   wire net_6884;
   wire net_6883;
   wire net_6882;
   wire net_6881;
   wire net_6880;
   wire net_6879;
   wire net_6878;
   wire net_6877;
   wire net_6876;
   wire net_6875;
   wire net_6874;
   wire net_6873;
   wire net_6872;
   wire net_6871;
   wire net_6870;
   wire net_6869;
   wire net_6868;
   wire net_6867;
   wire net_6866;
   wire net_6865;
   wire net_6864;
   wire net_6863;
   wire net_6862;
   wire net_6861;
   wire net_6860;
   wire net_6859;
   wire net_6858;
   wire net_6857;
   wire net_6856;
   wire net_6855;
   wire net_6854;
   wire net_6853;
   wire net_6852;
   wire net_6851;
   wire net_6850;
   wire net_6849;
   wire net_6848;
   wire net_6847;
   wire net_6846;
   wire net_6845;
   wire net_6844;
   wire net_6843;
   wire net_6842;
   wire net_6841;
   wire net_6840;
   wire net_6839;
   wire net_6838;
   wire net_6837;
   wire net_6836;
   wire net_6835;
   wire net_6834;
   wire net_6833;
   wire net_6832;
   wire net_6831;
   wire net_6830;
   wire net_6829;
   wire net_6826;
   wire net_6821;
   wire net_6820;
   wire net_6819;
   wire net_6818;
   wire net_6817;
   wire net_6816;
   wire net_6815;
   wire net_6814;
   wire net_6813;
   wire net_6812;
   wire net_6811;
   wire net_6810;
   wire net_6809;
   wire net_6808;
   wire net_6807;
   wire net_6806;
   wire net_6805;
   wire net_6804;
   wire net_6803;
   wire net_6802;
   wire net_6801;
   wire net_6800;
   wire net_6799;
   wire net_6798;
   wire net_6797;
   wire net_6796;
   wire net_6795;
   wire net_6794;
   wire net_6793;
   wire net_6792;
   wire net_6791;
   wire net_6790;
   wire net_6789;
   wire net_6788;
   wire net_6787;
   wire net_6786;
   wire net_6785;
   wire net_6784;
   wire net_6783;
   wire net_6782;
   wire net_6781;
   wire net_6780;
   wire net_6779;
   wire net_6778;
   wire net_6777;
   wire net_6776;
   wire net_6775;
   wire net_6774;
   wire net_6773;
   wire net_6772;
   wire net_6771;
   wire net_6770;
   wire net_6769;
   wire net_6768;
   wire net_6767;
   wire net_6766;
   wire net_6765;
   wire net_6764;
   wire net_6763;
   wire net_6762;
   wire net_6761;
   wire net_6760;
   wire net_6759;
   wire net_6758;
   wire net_6757;
   wire net_6756;
   wire net_6755;
   wire net_6754;
   wire net_6753;
   wire net_6752;
   wire net_6751;
   wire net_6750;
   wire net_6749;
   wire net_6748;
   wire net_6747;
   wire net_6746;
   wire net_6745;
   wire net_6744;
   wire net_6743;
   wire net_6742;
   wire net_6741;
   wire net_6740;
   wire net_6739;
   wire net_6738;
   wire net_6737;
   wire net_6736;
   wire net_6735;
   wire net_6734;
   wire net_6733;
   wire net_6732;
   wire net_6731;
   wire net_6730;
   wire net_6729;
   wire net_6728;
   wire net_6727;
   wire net_6726;
   wire net_6725;
   wire net_6724;
   wire net_6723;
   wire net_6722;
   wire net_6721;
   wire net_6720;
   wire net_6719;
   wire net_6718;
   wire net_6717;
   wire net_6716;
   wire net_6715;
   wire net_6714;
   wire net_6713;
   wire net_6712;
   wire net_6711;
   wire net_6710;
   wire net_6709;
   wire net_6708;
   wire net_6707;
   wire net_6706;
   wire net_6705;
   wire net_6704;
   wire net_6703;
   wire net_6702;
   wire net_6701;
   wire net_6700;
   wire net_6699;
   wire net_6698;
   wire net_6697;
   wire net_6696;
   wire net_6695;
   wire net_6694;
   wire net_6691;
   wire net_6686;
   wire net_6685;
   wire net_6684;
   wire net_6683;
   wire net_6682;
   wire net_6681;
   wire net_6680;
   wire net_6679;
   wire net_6678;
   wire net_6677;
   wire net_6676;
   wire net_6675;
   wire net_6674;
   wire net_6673;
   wire net_6672;
   wire net_6671;
   wire net_6670;
   wire net_6669;
   wire net_6668;
   wire net_6667;
   wire net_6666;
   wire net_6665;
   wire net_6664;
   wire net_6663;
   wire net_6662;
   wire net_6661;
   wire net_6660;
   wire net_6659;
   wire net_6658;
   wire net_6657;
   wire net_6656;
   wire net_6655;
   wire net_6654;
   wire net_6653;
   wire net_6652;
   wire net_6651;
   wire net_6650;
   wire net_6649;
   wire net_6648;
   wire net_6647;
   wire net_6646;
   wire net_6645;
   wire net_6644;
   wire net_6643;
   wire net_6642;
   wire net_6641;
   wire net_6640;
   wire net_6639;
   wire net_6638;
   wire net_6637;
   wire net_6636;
   wire net_6635;
   wire net_6634;
   wire net_6633;
   wire net_6632;
   wire net_6631;
   wire net_6630;
   wire net_6629;
   wire net_6628;
   wire net_6627;
   wire net_6626;
   wire net_6625;
   wire net_6624;
   wire net_6623;
   wire net_6622;
   wire net_6621;
   wire net_6620;
   wire net_6619;
   wire net_6618;
   wire net_6617;
   wire net_6616;
   wire net_6615;
   wire net_6614;
   wire net_6613;
   wire net_6612;
   wire net_6611;
   wire net_6610;
   wire net_6609;
   wire net_6608;
   wire net_6607;
   wire net_6606;
   wire net_6605;
   wire net_6604;
   wire net_6603;
   wire net_6602;
   wire net_6601;
   wire net_6600;
   wire net_6599;
   wire net_6598;
   wire net_6597;
   wire net_6596;
   wire net_6595;
   wire net_6594;
   wire net_6593;
   wire net_6592;
   wire net_6591;
   wire net_6590;
   wire net_6589;
   wire net_6588;
   wire net_6587;
   wire net_6586;
   wire net_6585;
   wire net_6584;
   wire net_6583;
   wire net_6582;
   wire net_6581;
   wire net_6580;
   wire net_6579;
   wire net_6578;
   wire net_6577;
   wire net_6576;
   wire net_6575;
   wire net_6574;
   wire net_6573;
   wire net_6572;
   wire net_6571;
   wire net_6570;
   wire net_6569;
   wire net_6568;
   wire net_6567;
   wire net_6566;
   wire net_6565;
   wire net_6564;
   wire net_6563;
   wire net_6562;
   wire net_6561;
   wire net_6560;
   wire net_6559;
   wire net_6556;
   wire net_6551;
   wire net_6550;
   wire net_6549;
   wire net_6548;
   wire net_6547;
   wire net_6546;
   wire net_6545;
   wire net_6544;
   wire net_6543;
   wire net_6542;
   wire net_6541;
   wire net_6540;
   wire net_6539;
   wire net_6538;
   wire net_6537;
   wire net_6536;
   wire net_6535;
   wire net_6534;
   wire net_6533;
   wire net_6532;
   wire net_6531;
   wire net_6530;
   wire net_6529;
   wire net_6528;
   wire net_6527;
   wire net_6526;
   wire net_6525;
   wire net_6524;
   wire net_6523;
   wire net_6522;
   wire net_6521;
   wire net_6520;
   wire net_6519;
   wire net_6518;
   wire net_6517;
   wire net_6516;
   wire net_6515;
   wire net_6514;
   wire net_6513;
   wire net_6512;
   wire net_6511;
   wire net_6510;
   wire net_6509;
   wire net_6508;
   wire net_6507;
   wire net_6506;
   wire net_6505;
   wire net_6504;
   wire net_6503;
   wire net_6502;
   wire net_6501;
   wire net_6500;
   wire net_6499;
   wire net_6498;
   wire net_6497;
   wire net_6496;
   wire net_6495;
   wire net_6494;
   wire net_6493;
   wire net_6492;
   wire net_6491;
   wire net_6490;
   wire net_6489;
   wire net_6488;
   wire net_6487;
   wire net_6486;
   wire net_6485;
   wire net_6484;
   wire net_6483;
   wire net_6482;
   wire net_6481;
   wire net_6480;
   wire net_6479;
   wire net_6478;
   wire net_6477;
   wire net_6476;
   wire net_6475;
   wire net_6474;
   wire net_6473;
   wire net_6472;
   wire net_6471;
   wire net_6470;
   wire net_6469;
   wire net_6468;
   wire net_6467;
   wire net_6466;
   wire net_6465;
   wire net_6464;
   wire net_6463;
   wire net_6462;
   wire net_6461;
   wire net_6460;
   wire net_6459;
   wire net_6458;
   wire net_6457;
   wire net_6456;
   wire net_6455;
   wire net_6454;
   wire net_6453;
   wire net_6452;
   wire net_6451;
   wire net_6450;
   wire net_6449;
   wire net_6448;
   wire net_6447;
   wire net_6446;
   wire net_6445;
   wire net_6444;
   wire net_6443;
   wire net_6442;
   wire net_6441;
   wire net_6440;
   wire net_6439;
   wire net_6438;
   wire net_6437;
   wire net_6436;
   wire net_6435;
   wire net_6434;
   wire net_6433;
   wire net_6432;
   wire net_6431;
   wire net_6430;
   wire net_6429;
   wire net_6428;
   wire net_6427;
   wire net_6426;
   wire net_6425;
   wire net_6424;
   wire net_6417;
   wire net_6416;
   wire net_6412;
   wire net_6403;
   wire net_6400;
   wire net_6399;
   wire net_6398;
   wire net_6397;
   wire net_6396;
   wire net_6395;
   wire net_6394;
   wire net_6393;
   wire net_6392;
   wire net_6391;
   wire net_6390;
   wire net_6389;
   wire net_6388;
   wire net_6387;
   wire net_6386;
   wire net_6385;
   wire net_6384;
   wire net_6383;
   wire net_6382;
   wire net_6381;
   wire net_6380;
   wire net_6379;
   wire net_6378;
   wire net_6377;
   wire net_6376;
   wire net_6375;
   wire net_6374;
   wire net_6373;
   wire net_6372;
   wire net_6371;
   wire net_6370;
   wire net_6369;
   wire net_6368;
   wire net_6367;
   wire net_6366;
   wire net_6365;
   wire net_6364;
   wire net_6363;
   wire net_6362;
   wire net_6361;
   wire net_6360;
   wire net_6359;
   wire net_6358;
   wire net_6357;
   wire net_6356;
   wire net_6355;
   wire net_6354;
   wire net_6353;
   wire net_6352;
   wire net_6351;
   wire net_6350;
   wire net_6349;
   wire net_6348;
   wire net_6347;
   wire net_6346;
   wire net_6345;
   wire net_6344;
   wire net_6343;
   wire net_6342;
   wire net_6341;
   wire net_6340;
   wire net_6339;
   wire net_6338;
   wire net_6337;
   wire net_6336;
   wire net_6335;
   wire net_6334;
   wire net_6333;
   wire net_6332;
   wire net_6331;
   wire net_6330;
   wire net_6329;
   wire net_6328;
   wire net_6327;
   wire net_6326;
   wire net_6325;
   wire net_6324;
   wire net_6323;
   wire net_6322;
   wire net_6321;
   wire net_6320;
   wire net_6318;
   wire net_6317;
   wire net_6316;
   wire net_6315;
   wire net_6314;
   wire net_6313;
   wire net_6312;
   wire net_6311;
   wire net_6310;
   wire net_6309;
   wire net_6308;
   wire net_6307;
   wire net_6306;
   wire net_6305;
   wire net_6304;
   wire net_6303;
   wire net_6302;
   wire net_6301;
   wire net_6300;
   wire net_6299;
   wire net_6279;
   wire net_6278;
   wire net_6277;
   wire net_6276;
   wire net_6275;
   wire net_6274;
   wire net_6273;
   wire net_6272;
   wire net_6271;
   wire net_6270;
   wire net_6269;
   wire net_6268;
   wire net_6267;
   wire net_6266;
   wire net_6265;
   wire net_6264;
   wire net_6263;
   wire net_6262;
   wire net_6261;
   wire net_6260;
   wire net_6258;
   wire net_6257;
   wire net_6256;
   wire net_6255;
   wire net_6254;
   wire net_6253;
   wire net_6252;
   wire net_6251;
   wire net_6250;
   wire net_6249;
   wire net_6248;
   wire net_6247;
   wire net_6246;
   wire net_6245;
   wire net_6244;
   wire net_6243;
   wire net_6242;
   wire net_6241;
   wire net_6240;
   wire net_6238;
   wire net_6237;
   wire net_6236;
   wire net_6235;
   wire net_6234;
   wire net_6233;
   wire net_6232;
   wire net_6231;
   wire net_6230;
   wire net_6229;
   wire net_6228;
   wire net_6227;
   wire net_6226;
   wire net_6225;
   wire net_6224;
   wire net_6223;
   wire net_6218;
   wire net_6217;
   wire net_6216;
   wire net_6215;
   wire net_6214;
   wire net_6213;
   wire net_6212;
   wire net_6211;
   wire net_6198;
   wire net_6197;
   wire net_6196;
   wire net_6195;
   wire net_6193;
   wire net_6192;
   wire net_6191;
   wire net_6190;
   wire net_6061;
   wire net_6060;
   wire net_6059;
   wire net_6058;
   wire net_6057;
   wire net_6056;
   wire net_6055;
   wire net_6054;
   wire net_6053;
   wire net_6047;
   wire net_6046;
   wire net_6036;
   wire net_6035;
   wire net_6025;
   wire net_6024;
   wire net_6014;
   wire net_6013;
   wire net_6003;
   wire net_5992;
   wire net_5861;
   wire net_5860;
   wire net_5858;
   wire net_5849;
   wire net_391;
   wire net_390;
   wire net_389;
   wire net_388;
   wire net_387;
   wire net_386;
   wire net_385;
   wire net_384;
   wire net_383;
   wire net_382;
   wire net_381;
   wire net_380;
   wire net_379;
   wire net_378;
   wire net_377;
   wire net_376;
   wire net_375;
   wire net_374;
   wire net_373;
   wire net_372;
   wire net_371;
   wire net_370;
   wire net_369;
   wire net_368;
   wire net_367;
   wire net_366;
   wire net_365;
   wire net_364;
   wire net_363;
   wire net_362;
   wire net_361;
   wire net_360;
   wire net_359;
   wire net_358;
   wire net_357;
   wire net_356;
   wire net_355;
   wire net_354;
   wire net_353;
   wire net_352;
   wire net_351;
   wire net_350;
   wire net_349;
   wire net_348;
   wire net_347;
   wire net_346;
   wire net_345;
   wire net_344;
   wire net_343;
   wire net_342;
   wire net_341;
   wire net_340;
   wire net_339;
   wire net_338;
   wire net_337;
   wire net_336;
   wire net_335;
   wire net_334;
   wire net_333;
   wire net_332;
   wire net_331;
   wire net_330;
   wire net_329;
   wire net_328;
   wire net_327;
   wire net_326;
   wire net_325;
   wire net_324;
   wire net_323;
   wire net_322;
   wire net_321;
   wire net_320;
   wire net_319;
   wire net_318;
   wire net_317;
   wire net_316;
   wire net_315;
   wire net_314;
   wire net_313;
   wire net_312;
   wire net_311;
   wire net_310;
   wire net_309;
   wire net_308;
   wire net_307;
   wire net_306;
   wire net_305;
   wire net_304;
   wire net_303;
   wire net_302;
   wire net_301;
   wire net_300;
   wire net_297;
   wire net_296;
   wire net_286;
   wire net_285;
   wire net_275;
   wire net_274;
   wire net_261;
   wire net_260;
   wire net_259;
   wire net_258;
   wire net_257;
   wire net_256;
   wire net_255;
   wire net_254;
   wire net_253;
   wire net_252;
   wire net_251;
   wire net_250;
   wire net_249;
   wire net_248;
   wire net_247;
   wire net_246;
   wire net_245;
   wire net_244;
   wire net_243;
   wire net_242;
   wire net_241;
   wire net_240;
   wire net_239;
   wire net_238;
   wire net_237;
   wire net_236;
   wire net_235;
   wire net_234;
   wire net_233;
   wire net_232;
   wire net_231;
   wire net_230;
   wire net_224;
   wire net_223;
   wire net_222;
   wire net_220;
   wire net_219;
   wire net_218;
   wire net_216;
   wire net_208;
   wire net_207;
   wire net_206;
   wire net_205;
   wire net_204;
   wire net_203;
   wire net_202;
   wire net_200;
   wire net_199;
   wire net_198;
   wire net_197;
   wire net_196;
   wire net_195;
   wire net_194;
   wire net_187;
   wire net_186;
   wire net_185;
   wire net_183;
   wire net_182;
   wire net_181;
   wire net_179;
   wire net_171;
   wire net_170;
   wire net_169;
   wire net_168;
   wire net_167;
   wire net_166;
   wire net_165;
   wire net_164;
   wire net_163;
   wire net_162;
   wire net_161;
   wire net_160;
   wire net_159;
   wire net_158;
   wire net_157;
   wire net_156;
   wire net_155;
   wire net_153;
   wire net_152;
   wire net_151;
   wire net_150;
   wire net_149;
   wire net_148;
   wire net_147;
   wire net_146;
   wire net_145;
   wire net_144;
   wire net_143;
   wire net_142;
   wire net_141;
   wire net_140;
   wire net_139;
   wire net_138;
   wire net_137;
   wire net_136;
   wire net_135;
   wire net_134;
   wire net_133;
   wire net_132;
   wire net_131;
   wire net_130;
   wire n9997;
   wire n9992;
   wire n9988;
   wire n9985;
   wire n9981;
   wire n9976;
   wire n9971;
   wire n9966;
   wire n9961;
   wire n9957;
   wire n9953;
   wire n995;
   wire n9949;
   wire n9944;
   wire n9939;
   wire n9935;
   wire n9930;
   wire n9926;
   wire n9923;
   wire n9918;
   wire n9914;
   wire n9911;
   wire n9907;
   wire n9902;
   wire n990;
   wire n9899;
   wire n9894;
   wire n9889;
   wire n9885;
   wire n9880;
   wire n9875;
   wire n9871;
   wire n9867;
   wire n9863;
   wire n9858;
   wire n9853;
   wire n985;
   wire n9849;
   wire n9844;
   wire n9840;
   wire n9837;
   wire n9833;
   wire n9828;
   wire n9824;
   wire n9819;
   wire n9814;
   wire n981;
   wire n9809;
   wire n9805;
   wire n9801;
   wire n9796;
   wire n9792;
   wire n9787;
   wire n9783;
   wire n9778;
   wire n9773;
   wire n9768;
   wire n9763;
   wire n976;
   wire n9758;
   wire n9754;
   wire n9750;
   wire n9746;
   wire n9742;
   wire n9737;
   wire n9733;
   wire n9729;
   wire n9724;
   wire n9719;
   wire n9714;
   wire n971;
   wire n9709;
   wire n9704;
   wire n9700;
   wire n9695;
   wire n9692;
   wire n9687;
   wire n9683;
   wire n9678;
   wire n9673;
   wire n9668;
   wire n9664;
   wire n9660;
   wire n966;
   wire n9655;
   wire n9651;
   wire n9647;
   wire n9642;
   wire n9638;
   wire n9633;
   wire n9628;
   wire n9624;
   wire n9620;
   wire n9616;
   wire n9611;
   wire n961;
   wire n9606;
   wire n9602;
   wire n9597;
   wire n9592;
   wire n9588;
   wire n9583;
   wire n9579;
   wire n9574;
   wire n9569;
   wire n9564;
   wire n956;
   wire n9559;
   wire n9554;
   wire n9549;
   wire n9546;
   wire n9541;
   wire n9537;
   wire n9533;
   wire n953;
   wire n9528;
   wire n9525;
   wire n9520;
   wire n9517;
   wire n9512;
   wire n9507;
   wire n9502;
   wire n9497;
   wire n9492;
   wire n9487;
   wire n9483;
   wire n948;
   wire n9478;
   wire n9475;
   wire n9470;
   wire n9467;
   wire n9462;
   wire n9459;
   wire n9454;
   wire n9449;
   wire n9445;
   wire n9441;
   wire n944;
   wire n9436;
   wire n9431;
   wire n9428;
   wire n9425;
   wire n9420;
   wire n9415;
   wire n9410;
   wire n9405;
   wire n9402;
   wire n940;
   wire n9398;
   wire n9393;
   wire n9390;
   wire n9385;
   wire n9381;
   wire n9377;
   wire n9373;
   wire n9370;
   wire n9365;
   wire n9361;
   wire n9356;
   wire n9352;
   wire n935;
   wire n9348;
   wire n9343;
   wire n9339;
   wire n9335;
   wire n9330;
   wire n9326;
   wire n9321;
   wire n9316;
   wire n9312;
   wire n9307;
   wire n9302;
   wire n930;
   wire n9298;
   wire n9294;
   wire n9290;
   wire n9287;
   wire n9282;
   wire n9277;
   wire n9272;
   wire n9267;
   wire n9263;
   wire n9258;
   wire n9254;
   wire n9250;
   wire n925;
   wire n9245;
   wire n9242;
   wire n9238;
   wire n9233;
   wire n9228;
   wire n9225;
   wire n9220;
   wire n9215;
   wire n9211;
   wire n9206;
   wire n9201;
   wire n920;
   wire n9196;
   wire n9192;
   wire n9187;
   wire n9182;
   wire n9178;
   wire n9173;
   wire n9169;
   wire n9164;
   wire n9160;
   wire n916;
   wire n9156;
   wire n9151;
   wire n9146;
   wire n9143;
   wire n9138;
   wire n9134;
   wire n9129;
   wire n9124;
   wire n9120;
   wire n9115;
   wire n9110;
   wire n911;
   wire n9106;
   wire n9101;
   wire n9096;
   wire n9091;
   wire n9086;
   wire n9082;
   wire n9079;
   wire n9074;
   wire n907;
   wire n9069;
   wire n9065;
   wire n9060;
   wire n9057;
   wire n9052;
   wire n9047;
   wire n9042;
   wire n9037;
   wire n9034;
   wire n9030;
   wire n903;
   wire n9025;
   wire n9022;
   wire n9017;
   wire n9014;
   wire n9010;
   wire n9005;
   wire n9000;
   wire n8995;
   wire n8990;
   wire n899;
   wire n8986;
   wire n8981;
   wire n8976;
   wire n8971;
   wire n8967;
   wire n8963;
   wire n8958;
   wire n8953;
   wire n8948;
   wire n8943;
   wire n894;
   wire n8939;
   wire n8934;
   wire n8931;
   wire n8926;
   wire n8922;
   wire n8917;
   wire n8912;
   wire n8908;
   wire n8903;
   wire n890;
   wire n8899;
   wire n8895;
   wire n8891;
   wire n8886;
   wire n8882;
   wire n8877;
   wire n8873;
   wire n8869;
   wire n8864;
   wire n8860;
   wire n8855;
   wire n8850;
   wire n885;
   wire n8845;
   wire n8840;
   wire n8835;
   wire n8831;
   wire n8826;
   wire n8823;
   wire n8818;
   wire n8813;
   wire n8809;
   wire n8805;
   wire n8800;
   wire n880;
   wire n8797;
   wire n8793;
   wire n8788;
   wire n8784;
   wire n8780;
   wire n8775;
   wire n8771;
   wire n8767;
   wire n8762;
   wire n8757;
   wire n8753;
   wire n875;
   wire n8748;
   wire n8743;
   wire n8739;
   wire n8734;
   wire n8730;
   wire n8725;
   wire n8720;
   wire n8715;
   wire n8711;
   wire n8708;
   wire n8703;
   wire n870;
   wire n8698;
   wire n8694;
   wire n8689;
   wire n8685;
   wire n8681;
   wire n8676;
   wire n8671;
   wire n867;
   wire n8666;
   wire n8662;
   wire n8658;
   wire n8654;
   wire n8650;
   wire n8645;
   wire n8641;
   wire n8637;
   wire n8632;
   wire n8628;
   wire n8625;
   wire n8621;
   wire n862;
   wire n8616;
   wire n8612;
   wire n8607;
   wire n8602;
   wire n8598;
   wire n8593;
   wire n8588;
   wire n8583;
   wire n8578;
   wire n8575;
   wire n8570;
   wire n857;
   wire n8565;
   wire n8561;
   wire n8557;
   wire n8552;
   wire n8549;
   wire n8544;
   wire n8540;
   wire n854;
   wire n8535;
   wire n8531;
   wire n8526;
   wire n8522;
   wire n8517;
   wire n8513;
   wire n8508;
   wire n8504;
   wire n8499;
   wire n8494;
   wire n8491;
   wire n849;
   wire n8486;
   wire n8481;
   wire n8477;
   wire n8472;
   wire n8467;
   wire n8464;
   wire n8459;
   wire n8455;
   wire n8451;
   wire n8447;
   wire n8443;
   wire n844;
   wire n8438;
   wire n8435;
   wire n8430;
   wire n8426;
   wire n8422;
   wire n8418;
   wire n8415;
   wire n8410;
   wire n8405;
   wire n8401;
   wire n8396;
   wire n8392;
   wire n839;
   wire n8387;
   wire n8382;
   wire n8377;
   wire n8372;
   wire n8367;
   wire n8362;
   wire n8359;
   wire n8354;
   wire n8350;
   wire n8345;
   wire n8340;
   wire n834;
   wire n8337;
   wire n8334;
   wire n8329;
   wire n8324;
   wire n8320;
   wire n8316;
   wire n8311;
   wire n8307;
   wire n8303;
   wire n830;
   wire n8299;
   wire n8294;
   wire n8289;
   wire n8284;
   wire n8280;
   wire n8276;
   wire n8271;
   wire n8266;
   wire n8262;
   wire n8258;
   wire n8253;
   wire n825;
   wire n8249;
   wire n8245;
   wire n8241;
   wire n8237;
   wire n8232;
   wire n8228;
   wire n8224;
   wire n8220;
   wire n8216;
   wire n8211;
   wire n8206;
   wire n8202;
   wire n820;
   wire n8197;
   wire n8192;
   wire n8188;
   wire n8183;
   wire n8179;
   wire n8174;
   wire n8170;
   wire n8166;
   wire n8161;
   wire n8156;
   wire n8152;
   wire n815;
   wire n8147;
   wire n8144;
   wire n8140;
   wire n8135;
   wire n8130;
   wire n8125;
   wire n8121;
   wire n8116;
   wire n8112;
   wire n811;
   wire n8107;
   wire n8102;
   wire n8097;
   wire n8092;
   wire n8088;
   wire n8085;
   wire n8080;
   wire n8075;
   wire n8072;
   wire n8067;
   wire n8064;
   wire n806;
   wire n8059;
   wire n8056;
   wire n8051;
   wire n8047;
   wire n8042;
   wire n8038;
   wire n8033;
   wire n8028;
   wire n8024;
   wire n802;
   wire n8019;
   wire n8015;
   wire n8010;
   wire n8005;
   wire n8002;
   wire n7997;
   wire n7994;
   wire n7989;
   wire n7985;
   wire n7980;
   wire n798;
   wire n7975;
   wire n7970;
   wire n7967;
   wire n7962;
   wire n7958;
   wire n7955;
   wire n7950;
   wire n7945;
   wire n7942;
   wire n7937;
   wire n7933;
   wire n793;
   wire n7929;
   wire n7924;
   wire n7920;
   wire n7916;
   wire n7911;
   wire n7906;
   wire n7902;
   wire n7897;
   wire n7893;
   wire n7888;
   wire n7883;
   wire n788;
   wire n7878;
   wire n7875;
   wire n7871;
   wire n7867;
   wire n7863;
   wire n7858;
   wire n7853;
   wire n7848;
   wire n7845;
   wire n7840;
   wire n7835;
   wire n7831;
   wire n783;
   wire n7826;
   wire n7822;
   wire n7818;
   wire n7815;
   wire n7810;
   wire n7806;
   wire n7802;
   wire n7798;
   wire n7793;
   wire n779;
   wire n7788;
   wire n7784;
   wire n7779;
   wire n7776;
   wire n7773;
   wire n7768;
   wire n7764;
   wire n7760;
   wire n7756;
   wire n7751;
   wire n7746;
   wire n7741;
   wire n774;
   wire n7737;
   wire n7732;
   wire n7728;
   wire n7723;
   wire n7719;
   wire n7714;
   wire n7709;
   wire n7704;
   wire n7700;
   wire n770;
   wire n7695;
   wire n7691;
   wire n7686;
   wire n7681;
   wire n7676;
   wire n7671;
   wire n7666;
   wire n7661;
   wire n7658;
   wire n7654;
   wire n765;
   wire n7649;
   wire n7644;
   wire n7640;
   wire n7635;
   wire n7631;
   wire n7626;
   wire n7622;
   wire n7618;
   wire n7613;
   wire n761;
   wire n7608;
   wire n7604;
   wire n7599;
   wire n7596;
   wire n7591;
   wire n7586;
   wire n7581;
   wire n7577;
   wire n7572;
   wire n7567;
   wire n7563;
   wire n756;
   wire n7558;
   wire n7553;
   wire n7548;
   wire n7543;
   wire n7539;
   wire n7535;
   wire n7530;
   wire n7527;
   wire n7522;
   wire n7518;
   wire n7513;
   wire n751;
   wire n7509;
   wire n7505;
   wire n7501;
   wire n7496;
   wire n7492;
   wire n7487;
   wire n7482;
   wire n7478;
   wire n7473;
   wire n7468;
   wire n7463;
   wire n746;
   wire n7459;
   wire n7454;
   wire n7450;
   wire n7446;
   wire n7442;
   wire n7437;
   wire n7432;
   wire n7427;
   wire n7422;
   wire n7417;
   wire n7413;
   wire n741;
   wire n7408;
   wire n7404;
   wire n7400;
   wire n7395;
   wire n7391;
   wire n7386;
   wire n7381;
   wire n7376;
   wire n7372;
   wire n7368;
   wire n7363;
   wire n736;
   wire n7359;
   wire n7354;
   wire n7349;
   wire n7344;
   wire n7340;
   wire n7335;
   wire n7330;
   wire n7326;
   wire n7321;
   wire n732;
   wire n7316;
   wire n7312;
   wire n7307;
   wire n7302;
   wire n7297;
   wire n7292;
   wire n7288;
   wire n7284;
   wire n7280;
   wire n7275;
   wire n7270;
   wire n727;
   wire n7265;
   wire n7260;
   wire n7256;
   wire n7252;
   wire n7249;
   wire n7245;
   wire n7240;
   wire n7235;
   wire n7230;
   wire n7226;
   wire n7221;
   wire n722;
   wire n7216;
   wire n7212;
   wire n7207;
   wire n7203;
   wire n7199;
   wire n7194;
   wire n7190;
   wire n7185;
   wire n7182;
   wire n718;
   wire n7177;
   wire n7172;
   wire n7167;
   wire n7164;
   wire n7160;
   wire n7155;
   wire n7151;
   wire n7147;
   wire n7142;
   wire n7138;
   wire n7133;
   wire n713;
   wire n7128;
   wire n7125;
   wire n7120;
   wire n7116;
   wire n7111;
   wire n7107;
   wire n7102;
   wire n7098;
   wire n7093;
   wire n7089;
   wire n7085;
   wire n7082;
   wire n708;
   wire n7077;
   wire n7072;
   wire n7067;
   wire n7062;
   wire n7058;
   wire n7053;
   wire n7049;
   wire n7045;
   wire n7041;
   wire n7036;
   wire n7032;
   wire n703;
   wire n7027;
   wire n7023;
   wire n7018;
   wire n7013;
   wire n7009;
   wire n7005;
   wire n7000;
   wire n6995;
   wire n6990;
   wire n6986;
   wire n6982;
   wire n698;
   wire n6977;
   wire n6974;
   wire n6969;
   wire n6964;
   wire n6960;
   wire n6957;
   wire n6952;
   wire n6947;
   wire n6943;
   wire n6938;
   wire n6934;
   wire n693;
   wire n6929;
   wire n6924;
   wire n6919;
   wire n6915;
   wire n6910;
   wire n6906;
   wire n6902;
   wire n6899;
   wire n6895;
   wire n6890;
   wire n6886;
   wire n6881;
   wire n688;
   wire n6876;
   wire n6872;
   wire n6867;
   wire n6863;
   wire n6860;
   wire n6855;
   wire n6850;
   wire n6845;
   wire n6840;
   wire n6836;
   wire n6831;
   wire n683;
   wire n6826;
   wire n6822;
   wire n6818;
   wire n6813;
   wire n6809;
   wire n6806;
   wire n6801;
   wire n6796;
   wire n6793;
   wire n6788;
   wire n6783;
   wire n678;
   wire n6779;
   wire n6774;
   wire n6770;
   wire n6765;
   wire n6761;
   wire n6756;
   wire n6752;
   wire n6749;
   wire n6746;
   wire n6741;
   wire n6736;
   wire n6732;
   wire n673;
   wire n6727;
   wire n6722;
   wire n6717;
   wire n6713;
   wire n6709;
   wire n6704;
   wire n6700;
   wire n6695;
   wire n6691;
   wire n669;
   wire n6687;
   wire n6682;
   wire n6678;
   wire n6674;
   wire n6669;
   wire n6665;
   wire n6661;
   wire n6656;
   wire n6652;
   wire n6648;
   wire n6643;
   wire n664;
   wire n6638;
   wire n6634;
   wire n6629;
   wire n6624;
   wire n6619;
   wire n6615;
   wire n6611;
   wire n6606;
   wire n6601;
   wire n6596;
   wire n6591;
   wire n659;
   wire n6586;
   wire n6583;
   wire n6578;
   wire n6574;
   wire n6570;
   wire n6566;
   wire n6563;
   wire n6558;
   wire n6554;
   wire n6550;
   wire n6545;
   wire n6540;
   wire n654;
   wire n6535;
   wire n6531;
   wire n6527;
   wire n6522;
   wire n6519;
   wire n6515;
   wire n6511;
   wire n6507;
   wire n6502;
   wire n6498;
   wire n6493;
   wire n649;
   wire n6489;
   wire n6485;
   wire n6480;
   wire n6477;
   wire n6472;
   wire n6469;
   wire n6464;
   wire n6460;
   wire n6455;
   wire n6450;
   wire n6446;
   wire n6441;
   wire n644;
   wire n6437;
   wire n6432;
   wire n6427;
   wire n6423;
   wire n6419;
   wire n6415;
   wire n6411;
   wire n6407;
   wire n6403;
   wire n6399;
   wire n6395;
   wire n6390;
   wire n639;
   wire n6386;
   wire n6381;
   wire n6376;
   wire n6371;
   wire n6367;
   wire n6362;
   wire n6357;
   wire n6354;
   wire n6350;
   wire n6346;
   wire n6342;
   wire n634;
   wire n6337;
   wire n6332;
   wire n6329;
   wire n6324;
   wire n6319;
   wire n6316;
   wire n6311;
   wire n6306;
   wire n6302;
   wire n6299;
   wire n6294;
   wire n6290;
   wire n629;
   wire n6285;
   wire n6281;
   wire n6276;
   wire n6271;
   wire n6266;
   wire n6261;
   wire n6258;
   wire n6254;
   wire n625;
   wire n6249;
   wire n6244;
   wire n6239;
   wire n6235;
   wire n6231;
   wire n6227;
   wire n6222;
   wire n6218;
   wire n6214;
   wire n6209;
   wire n6204;
   wire n6200;
   wire n620;
   wire n6195;
   wire n6191;
   wire n6186;
   wire n6181;
   wire n6176;
   wire n6171;
   wire n6166;
   wire n6161;
   wire n6158;
   wire n6153;
   wire n615;
   wire n6148;
   wire n6145;
   wire n6140;
   wire n6136;
   wire n6132;
   wire n6128;
   wire n6124;
   wire n6119;
   wire n6114;
   wire n6110;
   wire n6106;
   wire n6102;
   wire n610;
   wire n6098;
   wire n6093;
   wire n6088;
   wire n6083;
   wire n6078;
   wire n6074;
   wire n6069;
   wire n6066;
   wire n6061;
   wire n6056;
   wire n6052;
   wire n605;
   wire n6047;
   wire n6043;
   wire n6038;
   wire n6034;
   wire n6029;
   wire n6024;
   wire n6019;
   wire n6014;
   wire n6009;
   wire n6006;
   wire n6002;
   wire n600;
   wire n5997;
   wire n5992;
   wire n5987;
   wire n5982;
   wire n5978;
   wire n5973;
   wire n5968;
   wire n5964;
   wire n5960;
   wire n5955;
   wire n5951;
   wire n595;
   wire n5947;
   wire n5943;
   wire n5938;
   wire n5934;
   wire n5930;
   wire n5925;
   wire n5920;
   wire n5917;
   wire n5912;
   wire n5908;
   wire n5903;
   wire n590;
   wire n5899;
   wire n5894;
   wire n5890;
   wire n5885;
   wire n5881;
   wire n5876;
   wire n5872;
   wire n5867;
   wire n5864;
   wire n5860;
   wire n5855;
   wire n5850;
   wire n585;
   wire n5845;
   wire n5840;
   wire n5836;
   wire n5833;
   wire n5828;
   wire n5824;
   wire n5819;
   wire n5814;
   wire n5809;
   wire n5805;
   wire n5801;
   wire n580;
   wire n5796;
   wire n5792;
   wire n5787;
   wire n5783;
   wire n5779;
   wire n5775;
   wire n5771;
   wire n5767;
   wire n5763;
   wire n576;
   wire n5758;
   wire n5753;
   wire n5748;
   wire n5744;
   wire n5739;
   wire n5735;
   wire n5731;
   wire n5727;
   wire n5722;
   wire n5717;
   wire n5713;
   wire n571;
   wire n5709;
   wire n5704;
   wire n5700;
   wire n5696;
   wire n5691;
   wire n5686;
   wire n5682;
   wire n5679;
   wire n5674;
   wire n5669;
   wire n5664;
   wire n5660;
   wire n566;
   wire n5655;
   wire n5651;
   wire n5648;
   wire n5643;
   wire n5638;
   wire n5633;
   wire n5628;
   wire n5623;
   wire n5618;
   wire n5613;
   wire n5610;
   wire n561;
   wire n5606;
   wire n5601;
   wire n5596;
   wire n5591;
   wire n5588;
   wire n5584;
   wire n5579;
   wire n5575;
   wire n5570;
   wire n5565;
   wire n5560;
   wire n556;
   wire n5556;
   wire n5552;
   wire n5547;
   wire n5543;
   wire n5539;
   wire n5534;
   wire n553;
   wire n5529;
   wire n5525;
   wire n5521;
   wire n5517;
   wire n5513;
   wire n5508;
   wire n5504;
   wire n5500;
   wire n5495;
   wire n5490;
   wire n5486;
   wire n5481;
   wire n548;
   wire n5477;
   wire n5472;
   wire n5469;
   wire n5464;
   wire n5460;
   wire n5455;
   wire n5451;
   wire n5446;
   wire n5441;
   wire n5437;
   wire n5433;
   wire n543;
   wire n5429;
   wire n5424;
   wire n5420;
   wire n5415;
   wire n5411;
   wire n5406;
   wire n5402;
   wire n5397;
   wire n5393;
   wire n5388;
   wire n5383;
   wire n5380;
   wire n538;
   wire n5375;
   wire n5370;
   wire n5366;
   wire n5362;
   wire n5358;
   wire n5353;
   wire n5349;
   wire n5344;
   wire n5339;
   wire n5335;
   wire n5330;
   wire n533;
   wire n5326;
   wire n5321;
   wire n5316;
   wire n5312;
   wire n5307;
   wire n5302;
   wire n5298;
   wire n5293;
   wire n5288;
   wire n5284;
   wire n528;
   wire n5279;
   wire n5274;
   wire n5269;
   wire n5265;
   wire n5261;
   wire n5256;
   wire n5251;
   wire n5246;
   wire n5242;
   wire n5239;
   wire n5234;
   wire n5230;
   wire n523;
   wire n5225;
   wire n5221;
   wire n5217;
   wire n5212;
   wire n5207;
   wire n5202;
   wire n5198;
   wire n5193;
   wire n5189;
   wire n5186;
   wire n5181;
   wire n518;
   wire n5178;
   wire n5173;
   wire n5169;
   wire n5164;
   wire n5159;
   wire n5156;
   wire n5151;
   wire n5148;
   wire n5143;
   wire n5139;
   wire n5134;
   wire n5130;
   wire n513;
   wire n5126;
   wire n5121;
   wire n5117;
   wire n5112;
   wire n5107;
   wire n5103;
   wire n5098;
   wire n5094;
   wire n5090;
   wire n5085;
   wire n5080;
   wire n508;
   wire n5075;
   wire n5070;
   wire n5066;
   wire n5061;
   wire n5056;
   wire n5053;
   wire n5048;
   wire n5045;
   wire n5040;
   wire n5035;
   wire n5031;
   wire n503;
   wire n5027;
   wire n5023;
   wire n5018;
   wire n5013;
   wire n5008;
   wire n5005;
   wire n5001;
   wire n4996;
   wire n4992;
   wire n4987;
   wire n4983;
   wire n498;
   wire n4979;
   wire n4974;
   wire n4969;
   wire n4965;
   wire n4961;
   wire n4957;
   wire n4952;
   wire n4947;
   wire n4944;
   wire n4940;
   wire n4936;
   wire n4931;
   wire n493;
   wire n4927;
   wire n4922;
   wire n4917;
   wire n4913;
   wire n4908;
   wire n4904;
   wire n4899;
   wire n4895;
   wire n4890;
   wire n4886;
   wire n4881;
   wire n488;
   wire n4877;
   wire n4872;
   wire n4867;
   wire n4862;
   wire n4857;
   wire n4853;
   wire n4848;
   wire n4843;
   wire n484;
   wire n4838;
   wire n4834;
   wire n4831;
   wire n4827;
   wire n4822;
   wire n4818;
   wire n4814;
   wire n4809;
   wire n4805;
   wire n4800;
   wire n4795;
   wire n4791;
   wire n479;
   wire n4787;
   wire n4782;
   wire n4778;
   wire n4774;
   wire n4769;
   wire n4765;
   wire n4760;
   wire n4755;
   wire n4750;
   wire n4745;
   wire n4742;
   wire n474;
   wire n4737;
   wire n4732;
   wire n4727;
   wire n4722;
   wire n4717;
   wire n4713;
   wire n4708;
   wire n4703;
   wire n470;
   wire n4699;
   wire n4694;
   wire n4690;
   wire n4686;
   wire n4681;
   wire n4678;
   wire n4673;
   wire n4669;
   wire n4665;
   wire n4660;
   wire n4656;
   wire n4651;
   wire n465;
   wire n4646;
   wire n4641;
   wire n4636;
   wire n4631;
   wire n4627;
   wire n4622;
   wire n4617;
   wire n4613;
   wire n4609;
   wire n4604;
   wire n4600;
   wire n460;
   wire n4596;
   wire n4591;
   wire n4586;
   wire n4581;
   wire n4577;
   wire n4572;
   wire n4567;
   wire n4562;
   wire n4558;
   wire n4553;
   wire n455;
   wire n4548;
   wire n4544;
   wire n4539;
   wire n4534;
   wire n4529;
   wire n4524;
   wire n4520;
   wire n4515;
   wire n4510;
   wire n451;
   wire n4505;
   wire n4501;
   wire n4496;
   wire n4491;
   wire n4487;
   wire n4482;
   wire n4478;
   wire n4473;
   wire n447;
   wire n4469;
   wire n4464;
   wire n4459;
   wire n4456;
   wire n4451;
   wire n4448;
   wire n4443;
   wire n4438;
   wire n4433;
   wire n443;
   wire n4428;
   wire n4424;
   wire n4419;
   wire n4414;
   wire n4410;
   wire n4405;
   wire n4401;
   wire n4397;
   wire n4392;
   wire n4388;
   wire n4384;
   wire n438;
   wire n4379;
   wire n4374;
   wire n4370;
   wire n4365;
   wire n4362;
   wire n4357;
   wire n4352;
   wire n4348;
   wire n4343;
   wire n434;
   wire n4338;
   wire n4333;
   wire n4330;
   wire n4326;
   wire n4322;
   wire n4318;
   wire n4313;
   wire n4309;
   wire n4304;
   wire n4299;
   wire n4294;
   wire n429;
   wire n4289;
   wire n4284;
   wire n4280;
   wire n4276;
   wire n4271;
   wire n4267;
   wire n4263;
   wire n4258;
   wire n4253;
   wire n4249;
   wire n4245;
   wire n4240;
   wire n424;
   wire n4235;
   wire n4231;
   wire n4226;
   wire n4221;
   wire n4217;
   wire n4212;
   wire n4207;
   wire n4203;
   wire n420;
   wire n4199;
   wire n4194;
   wire n4191;
   wire n4186;
   wire n4181;
   wire n4176;
   wire n4171;
   wire n4166;
   wire n4161;
   wire n4158;
   wire n4153;
   wire n415;
   wire n4148;
   wire n4145;
   wire n4140;
   wire n4135;
   wire n4131;
   wire n4126;
   wire n4121;
   wire n4116;
   wire n4112;
   wire n4107;
   wire n4102;
   wire n410;
   wire n4098;
   wire n4094;
   wire n4089;
   wire n4084;
   wire n4079;
   wire n4075;
   wire n4071;
   wire n4068;
   wire n4063;
   wire n4059;
   wire n4055;
   wire n4051;
   wire n405;
   wire n4046;
   wire n4042;
   wire n4037;
   wire n4033;
   wire n4029;
   wire n4024;
   wire n4020;
   wire n4016;
   wire n4011;
   wire n4007;
   wire n4002;
   wire n400;
   wire n3998;
   wire n3993;
   wire n3989;
   wire n3985;
   wire n3981;
   wire n3976;
   wire n3972;
   wire n3967;
   wire n3962;
   wire n3957;
   wire n3953;
   wire n395;
   wire n3949;
   wire n3945;
   wire n3941;
   wire n3936;
   wire n3932;
   wire n3927;
   wire n3922;
   wire n3917;
   wire n3913;
   wire n3908;
   wire n3904;
   wire n390;
   wire n3899;
   wire n3896;
   wire n3891;
   wire n3886;
   wire n3881;
   wire n3877;
   wire n3872;
   wire n3867;
   wire n3864;
   wire n3859;
   wire n3855;
   wire n3851;
   wire n385;
   wire n3846;
   wire n3841;
   wire n3836;
   wire n3831;
   wire n3827;
   wire n3822;
   wire n3817;
   wire n3813;
   wire n3809;
   wire n3805;
   wire n3801;
   wire n380;
   wire n3796;
   wire n3791;
   wire n3787;
   wire n3782;
   wire n3777;
   wire n3773;
   wire n3770;
   wire n3765;
   wire n3761;
   wire n3756;
   wire n3752;
   wire n375;
   wire n3747;
   wire n3742;
   wire n3737;
   wire n3733;
   wire n3729;
   wire n3725;
   wire n3720;
   wire n3716;
   wire n3711;
   wire n3707;
   wire n3703;
   wire n370;
   wire n3698;
   wire n3693;
   wire n3689;
   wire n3684;
   wire n3679;
   wire n3675;
   wire n3670;
   wire n3666;
   wire n3661;
   wire n366;
   wire n3658;
   wire n3655;
   wire n3651;
   wire n3647;
   wire n3642;
   wire n3638;
   wire n3633;
   wire n3628;
   wire n3623;
   wire n3618;
   wire n3614;
   wire n361;
   wire n3609;
   wire n3604;
   wire n3600;
   wire n3595;
   wire n3590;
   wire n3587;
   wire n3582;
   wire n3577;
   wire n3572;
   wire n357;
   wire n3567;
   wire n3564;
   wire n3559;
   wire n3555;
   wire n3551;
   wire n3546;
   wire n3542;
   wire n3537;
   wire n3532;
   wire n3528;
   wire n3524;
   wire n3520;
   wire n352;
   wire n3516;
   wire n3511;
   wire n3507;
   wire n3502;
   wire n3497;
   wire n3494;
   wire n349;
   wire n3489;
   wire n3484;
   wire n3479;
   wire n3474;
   wire n3469;
   wire n3464;
   wire n3459;
   wire n3455;
   wire n3450;
   wire n3445;
   wire n3440;
   wire n344;
   wire n3436;
   wire n3431;
   wire n3427;
   wire n3422;
   wire n3418;
   wire n3413;
   wire n3408;
   wire n3404;
   wire n3400;
   wire n3395;
   wire n3390;
   wire n339;
   wire n3386;
   wire n3383;
   wire n3379;
   wire n3374;
   wire n3370;
   wire n3365;
   wire n3361;
   wire n3356;
   wire n3352;
   wire n3348;
   wire n3343;
   wire n334;
   wire n3338;
   wire n3333;
   wire n3330;
   wire n3325;
   wire n3322;
   wire n3318;
   wire n3313;
   wire n3308;
   wire n3303;
   wire n3299;
   wire n3294;
   wire n3290;
   wire n329;
   wire n3285;
   wire n3280;
   wire n3276;
   wire n3272;
   wire n3268;
   wire n3263;
   wire n3258;
   wire n3254;
   wire n3249;
   wire n3244;
   wire n3240;
   wire n324;
   wire n3235;
   wire n3231;
   wire n3226;
   wire n3222;
   wire n3217;
   wire n3212;
   wire n3207;
   wire n3203;
   wire n3199;
   wire n3194;
   wire n3190;
   wire n319;
   wire n3186;
   wire n3182;
   wire n3178;
   wire n3174;
   wire n3170;
   wire n3165;
   wire n3162;
   wire n3157;
   wire n3152;
   wire n3148;
   wire n3143;
   wire n314;
   wire n3139;
   wire n3134;
   wire n3130;
   wire n3126;
   wire n3121;
   wire n3117;
   wire n3114;
   wire n3110;
   wire n3105;
   wire n3102;
   wire n310;
   wire n3097;
   wire n3092;
   wire n3087;
   wire n3082;
   wire n3078;
   wire n3074;
   wire n3069;
   wire n3065;
   wire n3061;
   wire n3056;
   wire n3052;
   wire n305;
   wire n3047;
   wire n3042;
   wire n3037;
   wire n3033;
   wire n3030;
   wire n3025;
   wire n3020;
   wire n3015;
   wire n3010;
   wire n3005;
   wire n3000;
   wire n300;
   wire n2996;
   wire n2991;
   wire n2986;
   wire n2981;
   wire n2976;
   wire n2972;
   wire n2967;
   wire n2963;
   wire n2958;
   wire n2953;
   wire n295;
   wire n2948;
   wire n2944;
   wire n2939;
   wire n2935;
   wire n2930;
   wire n2926;
   wire n2922;
   wire n2918;
   wire n2913;
   wire n291;
   wire n2908;
   wire n2904;
   wire n2900;
   wire n2895;
   wire n2890;
   wire n2885;
   wire n2882;
   wire n2877;
   wire n2873;
   wire n2869;
   wire n2864;
   wire n2860;
   wire n286;
   wire n2855;
   wire n2850;
   wire n2845;
   wire n2840;
   wire n2836;
   wire n2831;
   wire n2827;
   wire n2823;
   wire n2819;
   wire n2814;
   wire n2810;
   wire n281;
   wire n2805;
   wire n2801;
   wire n2797;
   wire n2792;
   wire n2788;
   wire n2784;
   wire n2781;
   wire n2776;
   wire n2771;
   wire n2767;
   wire n2762;
   wire n276;
   wire n2758;
   wire n2753;
   wire n2748;
   wire n2745;
   wire n2741;
   wire n2737;
   wire n2732;
   wire n2727;
   wire n2723;
   wire n2718;
   wire n2713;
   wire n271;
   wire n2709;
   wire n2705;
   wire n2701;
   wire n2696;
   wire n2692;
   wire n2687;
   wire n2682;
   wire n2679;
   wire n2675;
   wire n2670;
   wire n2665;
   wire n2660;
   wire n266;
   wire n2656;
   wire n2651;
   wire n2647;
   wire n2642;
   wire n2637;
   wire n2632;
   wire n2627;
   wire n2622;
   wire n2618;
   wire n2615;
   wire n2610;
   wire n2605;
   wire n2601;
   wire n2597;
   wire n2594;
   wire n2590;
   wire n2585;
   wire n2580;
   wire n2575;
   wire n2570;
   wire n2566;
   wire n2561;
   wire n2556;
   wire n2552;
   wire n2547;
   wire n2543;
   wire n2539;
   wire n2534;
   wire n2529;
   wire n2524;
   wire n2519;
   wire n2515;
   wire n2510;
   wire n2505;
   wire n2500;
   wire n2496;
   wire n2493;
   wire n2488;
   wire n2484;
   wire n2479;
   wire n2474;
   wire n2470;
   wire n2465;
   wire n2462;
   wire n2457;
   wire n2452;
   wire n2448;
   wire n2444;
   wire n2440;
   wire n2435;
   wire n2430;
   wire n2426;
   wire n2422;
   wire n2417;
   wire n2414;
   wire n2409;
   wire n2404;
   wire n2399;
   wire n2395;
   wire n2391;
   wire n2386;
   wire n2381;
   wire n2377;
   wire n2373;
   wire n2370;
   wire n2365;
   wire n2360;
   wire n2355;
   wire n2350;
   wire n2347;
   wire n2342;
   wire n2338;
   wire n2334;
   wire n2329;
   wire n2324;
   wire n2321;
   wire n2316;
   wire n2312;
   wire n2307;
   wire n2303;
   wire n2298;
   wire n2293;
   wire n2288;
   wire n2284;
   wire n2280;
   wire n2275;
   wire n2270;
   wire n2265;
   wire n2260;
   wire n2256;
   wire n2251;
   wire n2247;
   wire n2242;
   wire n2237;
   wire n2232;
   wire n2227;
   wire n2222;
   wire n2218;
   wire n2213;
   wire n2208;
   wire n2203;
   wire n2199;
   wire n2194;
   wire n2189;
   wire n2186;
   wire n2181;
   wire n2177;
   wire n2172;
   wire n2167;
   wire n2162;
   wire n2157;
   wire n2152;
   wire n2149;
   wire n2144;
   wire n2140;
   wire n2136;
   wire n2132;
   wire n2127;
   wire n2122;
   wire n2119;
   wire n2115;
   wire n2111;
   wire n2106;
   wire n2102;
   wire n2098;
   wire n2093;
   wire n2088;
   wire n2084;
   wire n2079;
   wire n2074;
   wire n2070;
   wire n2065;
   wire n2060;
   wire n2055;
   wire n2051;
   wire n2046;
   wire n2041;
   wire n2036;
   wire n2031;
   wire n2026;
   wire n2021;
   wire n2016;
   wire n2011;
   wire n2007;
   wire n2002;
   wire n1998;
   wire n1993;
   wire n1988;
   wire n1983;
   wire n1978;
   wire n1973;
   wire n1969;
   wire n1964;
   wire n1959;
   wire n1954;
   wire n1950;
   wire n1945;
   wire n1941;
   wire n1936;
   wire n1932;
   wire n1927;
   wire n1922;
   wire n1918;
   wire n1913;
   wire n1908;
   wire n1903;
   wire n1898;
   wire n1893;
   wire n1888;
   wire n1883;
   wire n1878;
   wire n1874;
   wire n1869;
   wire n1865;
   wire n1860;
   wire n1855;
   wire n1851;
   wire n1846;
   wire n1841;
   wire n1836;
   wire n1832;
   wire n1827;
   wire n1822;
   wire n1817;
   wire n1812;
   wire n1807;
   wire n1802;
   wire n1797;
   wire n1792;
   wire n1787;
   wire n1782;
   wire n1779;
   wire n1775;
   wire n1770;
   wire n1765;
   wire n1761;
   wire n1756;
   wire n1752;
   wire n1747;
   wire n1742;
   wire n1737;
   wire n1732;
   wire n1727;
   wire n1722;
   wire n1718;
   wire n1714;
   wire n1709;
   wire n1704;
   wire n1701;
   wire n1696;
   wire n1691;
   wire n1686;
   wire n1681;
   wire n1677;
   wire n1673;
   wire n1668;
   wire n1663;
   wire n1658;
   wire n1653;
   wire n1649;
   wire n1644;
   wire n1639;
   wire n1634;
   wire n1629;
   wire n1624;
   wire n1619;
   wire n1615;
   wire n1610;
   wire n1605;
   wire n1600;
   wire n1596;
   wire n1591;
   wire n1587;
   wire n1582;
   wire n1577;
   wire n1572;
   wire n1568;
   wire n1564;
   wire n1560;
   wire n1555;
   wire n1551;
   wire n1546;
   wire n1542;
   wire n1538;
   wire n1533;
   wire n1528;
   wire n1524;
   wire n1519;
   wire n1515;
   wire n1510;
   wire n1506;
   wire n1501;
   wire n1496;
   wire n1491;
   wire n1487;
   wire n1482;
   wire n1478;
   wire n1474;
   wire n1469;
   wire n1465;
   wire n1460;
   wire n1455;
   wire n1451;
   wire n1446;
   wire n1442;
   wire n1438;
   wire n1433;
   wire n1428;
   wire n1423;
   wire n1419;
   wire n1414;
   wire n1410;
   wire n1405;
   wire n1400;
   wire n1396;
   wire n1391;
   wire n1386;
   wire n1383;
   wire n1378;
   wire n1373;
   wire n1368;
   wire n1363;
   wire n1359;
   wire n1355;
   wire n1350;
   wire n1345;
   wire n1340;
   wire n1335;
   wire n1331;
   wire n1326;
   wire n1322;
   wire n1318;
   wire n1314;
   wire n1309;
   wire n1305;
   wire n1300;
   wire n1295;
   wire n1291;
   wire n1287;
   wire n1282;
   wire n1277;
   wire n1272;
   wire n1267;
   wire n1262;
   wire n1258;
   wire n1253;
   wire n1248;
   wire n1244;
   wire n1240;
   wire n1236;
   wire n1232;
   wire n1228;
   wire n1224;
   wire n1219;
   wire n1214;
   wire n1210;
   wire n1205;
   wire n1200;
   wire n1195;
   wire n1191;
   wire n1187;
   wire n1183;
   wire n1178;
   wire n1173;
   wire n1168;
   wire n1163;
   wire n1158;
   wire n1153;
   wire n1148;
   wire n1144;
   wire n1140;
   wire n1135;
   wire n1130;
   wire n1125;
   wire n1121;
   wire n1116;
   wire n1111;
   wire n1106;
   wire n1102;
   wire n1097;
   wire n1093;
   wire n1089;
   wire n1085;
   wire n1081;
   wire n1077;
   wire n1072;
   wire n1067;
   wire n1062;
   wire n1058;
   wire n1053;
   wire n1049;
   wire n1044;
   wire n1039;
   wire n1034;
   wire n1029;
   wire n1024;
   wire n1020;
   wire n10158;
   wire n10154;
   wire n10150;
   wire n1015;
   wire n10145;
   wire n10141;
   wire n10137;
   wire n10132;
   wire n10128;
   wire n10124;
   wire n10120;
   wire n10116;
   wire n10112;
   wire n10107;
   wire n10103;
   wire n1010;
   wire n10099;
   wire n10094;
   wire n10089;
   wire n10084;
   wire n10079;
   wire n10074;
   wire n10070;
   wire n10066;
   wire n10061;
   wire n10056;
   wire n10052;
   wire n1005;
   wire n10047;
   wire n10042;
   wire n10037;
   wire n10032;
   wire n10028;
   wire n10023;
   wire n10019;
   wire n10014;
   wire n10010;
   wire n10006;
   wire n10001;
   wire n1000;
   wire _net_7824;
   wire _net_7823;
   wire _net_7822;
   wire _net_7821;
   wire _net_7820;
   wire _net_7819;
   wire _net_7818;
   wire _net_7817;
   wire _net_7816;
   wire _net_7815;
   wire _net_7814;
   wire _net_7813;
   wire _net_7812;
   wire _net_7811;
   wire _net_7810;
   wire _net_7809;
   wire _net_7808;
   wire _net_7806;
   wire _net_7805;
   wire _net_7804;
   wire _net_7803;
   wire _net_7801;
   wire _net_7800;
   wire _net_7798;
   wire _net_7797;
   wire _net_7796;
   wire _net_7795;
   wire _net_7794;
   wire _net_7793;
   wire _net_7791;
   wire _net_7789;
   wire _net_7788;
   wire _net_7787;
   wire _net_7786;
   wire _net_7785;
   wire _net_7784;
   wire _net_7783;
   wire _net_7782;
   wire _net_7781;
   wire _net_7768;
   wire _net_7765;
   wire _net_7763;
   wire _net_7761;
   wire _net_7759;
   wire _net_7757;
   wire _net_7755;
   wire _net_7753;
   wire _net_7751;
   wire _net_7749;
   wire _net_7748;
   wire _net_7747;
   wire _net_7746;
   wire _net_7745;
   wire _net_7736;
   wire _net_7735;
   wire _net_7734;
   wire _net_7733;
   wire _net_7732;
   wire _net_7731;
   wire _net_7730;
   wire _net_7729;
   wire _net_7728;
   wire _net_7727;
   wire _net_7726;
   wire _net_7725;
   wire _net_7724;
   wire _net_7723;
   wire _net_7722;
   wire _net_7721;
   wire _net_7720;
   wire _net_7719;
   wire _net_7718;
   wire _net_7717;
   wire _net_7716;
   wire _net_7707;
   wire _net_7706;
   wire _net_7705;
   wire _net_7704;
   wire _net_7703;
   wire _net_7702;
   wire _net_7701;
   wire _net_7700;
   wire _net_7699;
   wire _net_7698;
   wire _net_7697;
   wire _net_7696;
   wire _net_7695;
   wire _net_7694;
   wire _net_7693;
   wire _net_7692;
   wire _net_7690;
   wire _net_7689;
   wire _net_7688;
   wire _net_7687;
   wire _net_7686;
   wire _net_7685;
   wire _net_7684;
   wire _net_7683;
   wire _net_7682;
   wire _net_7681;
   wire _net_7667;
   wire _net_7666;
   wire _net_7665;
   wire _net_7664;
   wire _net_7663;
   wire _net_7662;
   wire _net_7661;
   wire _net_7660;
   wire _net_7659;
   wire _net_7658;
   wire _net_7657;
   wire _net_7656;
   wire _net_7655;
   wire _net_7654;
   wire _net_7653;
   wire _net_7652;
   wire _net_7651;
   wire _net_7650;
   wire _net_7649;
   wire _net_7648;
   wire _net_7635;
   wire _net_7634;
   wire _net_7633;
   wire _net_7632;
   wire _net_7631;
   wire _net_7630;
   wire _net_7629;
   wire _net_7628;
   wire _net_7627;
   wire _net_7626;
   wire _net_7625;
   wire _net_7624;
   wire _net_7623;
   wire _net_7622;
   wire _net_7621;
   wire _net_7620;
   wire _net_7619;
   wire _net_7618;
   wire _net_7617;
   wire _net_7616;
   wire _net_7603;
   wire _net_7602;
   wire _net_7601;
   wire _net_7600;
   wire _net_7599;
   wire _net_7598;
   wire _net_7597;
   wire _net_7596;
   wire _net_7595;
   wire _net_7594;
   wire _net_7593;
   wire _net_7592;
   wire _net_7591;
   wire _net_7590;
   wire _net_7589;
   wire _net_7588;
   wire _net_7587;
   wire _net_7586;
   wire _net_7585;
   wire _net_7584;
   wire _net_7583;
   wire _net_7582;
   wire _net_7581;
   wire _net_7580;
   wire _net_7579;
   wire _net_7578;
   wire _net_7577;
   wire _net_7576;
   wire _net_7575;
   wire _net_7574;
   wire _net_7573;
   wire _net_7572;
   wire _net_7571;
   wire _net_7570;
   wire _net_7569;
   wire _net_7568;
   wire _net_7567;
   wire _net_7566;
   wire _net_7565;
   wire _net_7564;
   wire _net_7563;
   wire _net_7562;
   wire _net_7561;
   wire _net_7560;
   wire _net_7559;
   wire _net_7558;
   wire _net_7557;
   wire _net_7556;
   wire _net_7555;
   wire _net_7554;
   wire _net_7553;
   wire _net_7552;
   wire _net_7535;
   wire _net_7534;
   wire _net_7533;
   wire _net_7532;
   wire _net_7531;
   wire _net_7530;
   wire _net_7516;
   wire _net_7515;
   wire _net_7514;
   wire _net_7513;
   wire _net_7512;
   wire _net_7511;
   wire _net_7510;
   wire _net_7509;
   wire _net_7508;
   wire _net_7507;
   wire _net_7506;
   wire _net_7505;
   wire _net_7504;
   wire _net_7503;
   wire _net_7502;
   wire _net_7501;
   wire _net_7500;
   wire _net_7499;
   wire _net_7498;
   wire _net_7497;
   wire _net_7484;
   wire _net_7483;
   wire _net_7482;
   wire _net_7481;
   wire _net_7480;
   wire _net_7479;
   wire _net_7478;
   wire _net_7477;
   wire _net_7476;
   wire _net_7475;
   wire _net_7474;
   wire _net_7473;
   wire _net_7472;
   wire _net_7471;
   wire _net_7470;
   wire _net_7469;
   wire _net_7468;
   wire _net_7467;
   wire _net_7466;
   wire _net_7465;
   wire _net_7452;
   wire _net_7451;
   wire _net_7450;
   wire _net_7449;
   wire _net_7448;
   wire _net_7447;
   wire _net_7446;
   wire _net_7445;
   wire _net_7444;
   wire _net_7443;
   wire _net_7442;
   wire _net_7441;
   wire _net_7440;
   wire _net_7439;
   wire _net_7438;
   wire _net_7437;
   wire _net_7436;
   wire _net_7435;
   wire _net_7434;
   wire _net_7433;
   wire _net_7432;
   wire _net_7431;
   wire _net_7430;
   wire _net_7429;
   wire _net_7428;
   wire _net_7427;
   wire _net_7426;
   wire _net_7425;
   wire _net_7424;
   wire _net_7423;
   wire _net_7422;
   wire _net_7421;
   wire _net_7420;
   wire _net_7419;
   wire _net_7418;
   wire _net_7417;
   wire _net_7416;
   wire _net_7415;
   wire _net_7414;
   wire _net_7413;
   wire _net_7412;
   wire _net_7411;
   wire _net_7410;
   wire _net_7409;
   wire _net_7408;
   wire _net_7407;
   wire _net_7406;
   wire _net_7405;
   wire _net_7404;
   wire _net_7403;
   wire _net_7402;
   wire _net_7401;
   wire _net_7384;
   wire _net_7383;
   wire _net_7382;
   wire _net_7381;
   wire _net_7380;
   wire _net_7379;
   wire _net_7365;
   wire _net_7364;
   wire _net_7363;
   wire _net_7362;
   wire _net_7361;
   wire _net_7360;
   wire _net_7359;
   wire _net_7358;
   wire _net_7357;
   wire _net_7356;
   wire _net_7355;
   wire _net_7354;
   wire _net_7353;
   wire _net_7352;
   wire _net_7351;
   wire _net_7350;
   wire _net_7349;
   wire _net_7348;
   wire _net_7347;
   wire _net_7346;
   wire _net_7333;
   wire _net_7332;
   wire _net_7331;
   wire _net_7330;
   wire _net_7329;
   wire _net_7328;
   wire _net_7327;
   wire _net_7326;
   wire _net_7325;
   wire _net_7324;
   wire _net_7323;
   wire _net_7322;
   wire _net_7321;
   wire _net_7320;
   wire _net_7319;
   wire _net_7318;
   wire _net_7317;
   wire _net_7316;
   wire _net_7315;
   wire _net_7314;
   wire _net_7301;
   wire _net_7300;
   wire _net_7299;
   wire _net_7298;
   wire _net_7297;
   wire _net_7296;
   wire _net_7295;
   wire _net_7294;
   wire _net_7293;
   wire _net_7292;
   wire _net_7291;
   wire _net_7290;
   wire _net_7289;
   wire _net_7288;
   wire _net_7287;
   wire _net_7286;
   wire _net_7285;
   wire _net_7284;
   wire _net_7283;
   wire _net_7282;
   wire _net_7281;
   wire _net_7280;
   wire _net_7279;
   wire _net_7278;
   wire _net_7277;
   wire _net_7276;
   wire _net_7275;
   wire _net_7274;
   wire _net_7273;
   wire _net_7272;
   wire _net_7271;
   wire _net_7270;
   wire _net_7269;
   wire _net_7268;
   wire _net_7267;
   wire _net_7266;
   wire _net_7265;
   wire _net_7264;
   wire _net_7263;
   wire _net_7262;
   wire _net_7261;
   wire _net_7260;
   wire _net_7259;
   wire _net_7258;
   wire _net_7257;
   wire _net_7256;
   wire _net_7255;
   wire _net_7254;
   wire _net_7253;
   wire _net_7252;
   wire _net_7251;
   wire _net_7250;
   wire _net_7233;
   wire _net_7232;
   wire _net_7230;
   wire _net_7229;
   wire _net_7228;
   wire _net_7227;
   wire _net_7098;
   wire _net_7097;
   wire _net_7095;
   wire _net_7094;
   wire _net_7093;
   wire _net_7092;
   wire _net_6963;
   wire _net_6962;
   wire _net_6960;
   wire _net_6959;
   wire _net_6958;
   wire _net_6957;
   wire _net_6828;
   wire _net_6827;
   wire _net_6825;
   wire _net_6824;
   wire _net_6823;
   wire _net_6822;
   wire _net_6693;
   wire _net_6692;
   wire _net_6690;
   wire _net_6689;
   wire _net_6688;
   wire _net_6687;
   wire _net_6558;
   wire _net_6557;
   wire _net_6555;
   wire _net_6554;
   wire _net_6553;
   wire _net_6552;
   wire _net_6423;
   wire _net_6422;
   wire _net_6421;
   wire _net_6420;
   wire _net_6419;
   wire _net_6418;
   wire _net_6415;
   wire _net_6414;
   wire _net_6413;
   wire _net_6411;
   wire _net_6410;
   wire _net_6409;
   wire _net_6408;
   wire _net_6407;
   wire _net_6406;
   wire _net_6405;
   wire _net_6404;
   wire _net_6402;
   wire _net_6401;
   wire _net_6319;
   wire _net_6298;
   wire _net_6297;
   wire _net_6296;
   wire _net_6295;
   wire _net_6294;
   wire _net_6293;
   wire _net_6292;
   wire _net_6291;
   wire _net_6290;
   wire _net_6289;
   wire _net_6288;
   wire _net_6287;
   wire _net_6286;
   wire _net_6285;
   wire _net_6284;
   wire _net_6283;
   wire _net_6282;
   wire _net_6281;
   wire _net_6280;
   wire _net_6259;
   wire _net_6239;
   wire _net_6222;
   wire _net_6221;
   wire _net_6220;
   wire _net_6219;
   wire _net_6210;
   wire _net_6209;
   wire _net_6208;
   wire _net_6207;
   wire _net_6206;
   wire _net_6205;
   wire _net_6204;
   wire _net_6203;
   wire _net_6202;
   wire _net_6201;
   wire _net_6200;
   wire _net_6199;
   wire _net_6194;
   wire _net_6189;
   wire _net_6188;
   wire _net_6187;
   wire _net_6186;
   wire _net_6185;
   wire _net_6184;
   wire _net_6183;
   wire _net_6182;
   wire _net_6181;
   wire _net_6180;
   wire _net_6179;
   wire _net_6178;
   wire _net_6177;
   wire _net_6176;
   wire _net_6175;
   wire _net_6174;
   wire _net_6173;
   wire _net_6172;
   wire _net_6171;
   wire _net_6170;
   wire _net_6169;
   wire _net_6168;
   wire _net_6167;
   wire _net_6166;
   wire _net_6165;
   wire _net_6164;
   wire _net_6163;
   wire _net_6162;
   wire _net_6161;
   wire _net_6160;
   wire _net_6159;
   wire _net_6158;
   wire _net_6157;
   wire _net_6156;
   wire _net_6155;
   wire _net_6154;
   wire _net_6153;
   wire _net_6152;
   wire _net_6151;
   wire _net_6150;
   wire _net_6149;
   wire _net_6148;
   wire _net_6147;
   wire _net_6146;
   wire _net_6145;
   wire _net_6144;
   wire _net_6143;
   wire _net_6142;
   wire _net_6141;
   wire _net_6140;
   wire _net_6139;
   wire _net_6138;
   wire _net_6137;
   wire _net_6136;
   wire _net_6135;
   wire _net_6134;
   wire _net_6133;
   wire _net_6132;
   wire _net_6131;
   wire _net_6130;
   wire _net_6129;
   wire _net_6128;
   wire _net_6127;
   wire _net_6126;
   wire _net_6125;
   wire _net_6124;
   wire _net_6123;
   wire _net_6122;
   wire _net_6121;
   wire _net_6120;
   wire _net_6119;
   wire _net_6118;
   wire _net_6117;
   wire _net_6116;
   wire _net_6115;
   wire _net_6114;
   wire _net_6113;
   wire _net_6112;
   wire _net_6111;
   wire _net_6110;
   wire _net_6109;
   wire _net_6108;
   wire _net_6107;
   wire _net_6106;
   wire _net_6105;
   wire _net_6104;
   wire _net_6103;
   wire _net_6102;
   wire _net_6101;
   wire _net_6100;
   wire _net_6099;
   wire _net_6098;
   wire _net_6097;
   wire _net_6096;
   wire _net_6095;
   wire _net_6094;
   wire _net_6093;
   wire _net_6092;
   wire _net_6091;
   wire _net_6090;
   wire _net_6089;
   wire _net_6088;
   wire _net_6087;
   wire _net_6086;
   wire _net_6085;
   wire _net_6084;
   wire _net_6083;
   wire _net_6082;
   wire _net_6081;
   wire _net_6080;
   wire _net_6079;
   wire _net_6078;
   wire _net_6077;
   wire _net_6076;
   wire _net_6075;
   wire _net_6074;
   wire _net_6073;
   wire _net_6072;
   wire _net_6071;
   wire _net_6070;
   wire _net_6069;
   wire _net_6068;
   wire _net_6067;
   wire _net_6066;
   wire _net_6065;
   wire _net_6064;
   wire _net_6063;
   wire _net_6062;
   wire _net_6052;
   wire _net_6051;
   wire _net_6050;
   wire _net_6049;
   wire _net_6048;
   wire _net_6045;
   wire _net_6044;
   wire _net_6043;
   wire _net_6042;
   wire _net_6041;
   wire _net_6040;
   wire _net_6039;
   wire _net_6038;
   wire _net_6037;
   wire _net_6034;
   wire _net_6033;
   wire _net_6032;
   wire _net_6031;
   wire _net_6030;
   wire _net_6029;
   wire _net_6028;
   wire _net_6027;
   wire _net_6026;
   wire _net_6023;
   wire _net_6022;
   wire _net_6021;
   wire _net_6020;
   wire _net_6019;
   wire _net_6018;
   wire _net_6017;
   wire _net_6016;
   wire _net_6015;
   wire _net_6012;
   wire _net_6011;
   wire _net_6010;
   wire _net_6009;
   wire _net_6008;
   wire _net_6007;
   wire _net_6006;
   wire _net_6005;
   wire _net_6004;
   wire _net_6002;
   wire _net_6001;
   wire _net_6000;
   wire _net_5999;
   wire _net_5998;
   wire _net_5997;
   wire _net_5996;
   wire _net_5995;
   wire _net_5994;
   wire _net_5993;
   wire _net_5991;
   wire _net_5990;
   wire _net_5989;
   wire _net_5988;
   wire _net_5987;
   wire _net_5986;
   wire _net_5985;
   wire _net_5984;
   wire _net_5983;
   wire _net_5982;
   wire _net_5981;
   wire _net_5980;
   wire _net_5979;
   wire _net_5978;
   wire _net_5977;
   wire _net_5976;
   wire _net_5975;
   wire _net_5974;
   wire _net_5973;
   wire _net_5972;
   wire _net_5971;
   wire _net_5970;
   wire _net_5969;
   wire _net_5968;
   wire _net_5967;
   wire _net_5966;
   wire _net_5965;
   wire _net_5964;
   wire _net_5963;
   wire _net_5962;
   wire _net_5961;
   wire _net_5960;
   wire _net_5924;
   wire _net_5922;
   wire _net_5920;
   wire _net_5859;
   wire _net_5857;
   wire _net_5856;
   wire _net_5855;
   wire _net_5854;
   wire _net_5853;
   wire _net_5852;
   wire _net_5851;
   wire _net_5850;
   wire _net_5848;
   wire _net_392;
   wire _net_299;
   wire _net_298;
   wire _net_295;
   wire _net_294;
   wire _net_293;
   wire _net_292;
   wire _net_291;
   wire _net_290;
   wire _net_289;
   wire _net_288;
   wire _net_287;
   wire _net_284;
   wire _net_283;
   wire _net_282;
   wire _net_281;
   wire _net_280;
   wire _net_279;
   wire _net_278;
   wire _net_277;
   wire _net_276;
   wire _net_273;
   wire _net_272;
   wire _net_271;
   wire _net_270;
   wire _net_269;
   wire _net_268;
   wire _net_267;
   wire _net_266;
   wire _net_265;
   wire _net_264;
   wire _net_263;
   wire _net_262;
   wire _net_229;
   wire _net_228;
   wire _net_227;
   wire _net_226;
   wire _net_225;
   wire _net_221;
   wire _net_217;
   wire _net_215;
   wire _net_214;
   wire _net_213;
   wire _net_212;
   wire _net_211;
   wire _net_210;
   wire _net_209;
   wire _net_201;
   wire _net_193;
   wire _net_192;
   wire _net_191;
   wire _net_190;
   wire _net_189;
   wire _net_188;
   wire _net_184;
   wire _net_180;
   wire _net_178;
   wire _net_177;
   wire _net_176;
   wire _net_175;
   wire _net_174;
   wire _net_173;
   wire _net_172;
   wire _net_154;
   wire _net_129;
   wire _net_128;
   wire _net_127;
   wire _net_126;
   wire _net_125;
   wire _net_124;
   wire _net_123;
   wire _net_122;
   wire _net_121;
   wire _net_120;
   wire _net_119;
   wire _net_118;
   wire _net_117;
   wire _net_116;
   wire _net_115;
   wire _net_114;
   wire _net_113;
   wire ck_net_4_19_a_2;
   wire ck_net_4_19_b_1;
   wire ck_net_4_15_a_2;
   wire ck_net_4_22_b_1;
   wire ck_net_4_20_b_1;
   wire ck_net_4_15_b_1;
   wire ck_net_4_21_b_1;
   wire ck_net_4_18_b_1;
   wire ck_net_4_18_a_1;
   wire ck_net_4_17_b_1;
   wire ck_net_4_17_a_1;
   wire ck_net_4_16_b_1;
   wire ck_net_4_16_a_1;
   wire ck_net_4_14_a_2;
   wire ck_net_4_10_b_1;
   wire ck_net_4_14_b_1;
   wire ck_net_4_11_b_1;
   wire ck_net_4_12_a_2;
   wire ck_net_4_9_b_1;
   wire ck_net_4_7_b_1;
   wire ck_net_4_7_a_1;
   wire ck_net_4_13_b_1;
   wire ck_net_4_12_b_1;
   wire ck_net_4_8_b_1;
   wire ck_net_1_0_b_2;
   wire ck_net_1_0_a_2;
   wire ck_net_1_0_0;
   wire clk;

   // Assignments 

   // Module instantiations
   LOGIC1_X1 t0 (
	   .Z (n7265) );
   DFF_X1 l2199 (
	   .Q (net_7041),
	   .D (n10158),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2198 (
	   .Q (net_6772),
	   .D (n10154),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2197 (
	   .Q (_net_6164),
	   .D (n10150),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2196 (
	   .Q (net_7313),
	   .D (n10145),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l2195 (
	   .Q (_net_7793),
	   .D (n10141),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l2194 (
	   .Q (_net_6176),
	   .D (n10137),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l2193 (
	   .Q (net_6532),
	   .D (n10132),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l2192 (
	   .Q (_net_7356),
	   .D (n10128),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2191 (
	   .Q (net_148),
	   .D (n10124),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l2190 (
	   .Q (net_6780),
	   .D (n10120),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2189 (
	   .Q (net_248),
	   .D (n10116),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l2188 (
	   .Q (net_7112),
	   .D (n10112),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2187 (
	   .Q (net_6648),
	   .D (n10107),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l2186 (
	   .Q (net_6645),
	   .D (n10103),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l2185 (
	   .Q (_net_7479),
	   .D (n10099),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l2184 (
	   .Q (_net_7264),
	   .D (n10094),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2183 (
	   .Q (_net_6183),
	   .D (n10089),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l2182 (
	   .Q (_net_6131),
	   .D (n10084),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l2181 (
	   .Q (_net_6555),
	   .D (n10079),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l2180 (
	   .Q (_net_7251),
	   .D (n10074),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2179 (
	   .Q (net_6884),
	   .D (n10070),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l2178 (
	   .Q (x620),
	   .D (n10066),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l2177 (
	   .Q (net_7773),
	   .D (n10061),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l2176 (
	   .Q (net_7677),
	   .D (n10056),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l2175 (
	   .Q (_net_7287),
	   .D (n10052),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2174 (
	   .Q (net_6351),
	   .D (n10047),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l2173 (
	   .Q (_net_6203),
	   .D (n10042),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l2172 (
	   .Q (_net_6017),
	   .D (n10037),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l2171 (
	   .Q (_net_7582),
	   .D (n10032),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2170 (
	   .Q (net_6879),
	   .D (n10028),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l2169 (
	   .Q (net_6224),
	   .D (n10023),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l2168 (
	   .Q (_net_267),
	   .D (n10019),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l2167 (
	   .Q (_net_7823),
	   .D (n10014),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l2166 (
	   .Q (net_6529),
	   .D (n10010),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l2165 (
	   .Q (net_6198),
	   .D (n10006),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2164 (
	   .Q (net_6507),
	   .D (n10001),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l2163 (
	   .Q (_net_7717),
	   .D (n9997),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l2162 (
	   .Q (net_7175),
	   .D (n9992),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2161 (
	   .Q (net_6905),
	   .D (n9988),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l2160 (
	   .Q (net_6381),
	   .D (n9985),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l2159 (
	   .Q (_net_7788),
	   .D (n9981),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l2158 (
	   .Q (net_6192),
	   .D (n9976),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2157 (
	   .Q (_net_6076),
	   .D (n9971),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l2156 (
	   .Q (_net_7402),
	   .D (n9966),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l2155 (
	   .Q (net_7071),
	   .D (n9961),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l2154 (
	   .Q (net_354),
	   .D (n9957),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l2153 (
	   .Q (net_7740),
	   .D (n9953),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l2152 (
	   .Q (_net_7348),
	   .D (n9949),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2151 (
	   .Q (net_6370),
	   .D (n9944),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l2150 (
	   .Q (_net_288),
	   .D (n9939),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l2149 (
	   .Q (net_6465),
	   .D (n9935),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l2148 (
	   .Q (net_338),
	   .D (n9930),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2147 (
	   .Q (net_374),
	   .D (n9926),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l2146 (
	   .Q (net_6719),
	   .D (n9923),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2145 (
	   .Q (_net_7795),
	   .D (n9918),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l2144 (
	   .Q (net_7221),
	   .D (n9914),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l2143 (
	   .Q (net_6446),
	   .D (n9911),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l2142 (
	   .Q (x361),
	   .D (n9907),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2141 (
	   .Q (net_6795),
	   .D (n9902),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l2140 (
	   .Q (net_6752),
	   .D (n9899),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2139 (
	   .Q (_net_287),
	   .D (n9894),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l2138 (
	   .Q (_net_6111),
	   .D (n9889),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l2137 (
	   .Q (net_7109),
	   .D (n9885),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2136 (
	   .Q (_net_6421),
	   .D (n9880),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2135 (
	   .Q (net_6533),
	   .D (n9875),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2134 (
	   .Q (net_6929),
	   .D (n9871),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l2133 (
	   .Q (net_6943),
	   .D (n9867),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l2132 (
	   .Q (_net_7097),
	   .D (n9863),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2131 (
	   .Q (_net_6407),
	   .D (n9858),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l2130 (
	   .Q (net_7644),
	   .D (n9853),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2129 (
	   .Q (_net_7421),
	   .D (n9849),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l2128 (
	   .Q (net_305),
	   .D (n9844),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2127 (
	   .Q (net_321),
	   .D (n9840),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l2126 (
	   .Q (net_7122),
	   .D (n9837),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l2125 (
	   .Q (net_7135),
	   .D (n9833),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l2124 (
	   .Q (net_7674),
	   .D (n9828),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l2123 (
	   .Q (_net_7383),
	   .D (n9824),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l2122 (
	   .Q (_net_7533),
	   .D (n9819),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l2121 (
	   .Q (_net_5859),
	   .D (n9814),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l2120 (
	   .Q (net_313),
	   .D (n9809),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2119 (
	   .Q (net_384),
	   .D (n9805),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2118 (
	   .Q (_net_7384),
	   .D (n9801),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l2117 (
	   .Q (net_6807),
	   .D (n9796),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l2116 (
	   .Q (_net_5989),
	   .D (n9792),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l2115 (
	   .Q (_net_7566),
	   .D (n9787),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l2114 (
	   .Q (net_7027),
	   .D (n9783),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l2113 (
	   .Q (_net_5973),
	   .D (n9778),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l2112 (
	   .Q (_net_6002),
	   .D (n9773),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l2111 (
	   .Q (_net_7283),
	   .D (n9768),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2110 (
	   .Q (_net_7576),
	   .D (n9763),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l2109 (
	   .Q (net_7669),
	   .D (n9758),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l2108 (
	   .Q (net_7522),
	   .D (n9754),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l2107 (
	   .Q (net_6657),
	   .D (n9750),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l2106 (
	   .Q (net_7214),
	   .D (n9746),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l2105 (
	   .Q (net_170),
	   .D (n9742),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2104 (
	   .Q (_net_7817),
	   .D (n9737),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l2103 (
	   .Q (_net_192),
	   .D (n9733),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l2102 (
	   .Q (net_6472),
	   .D (n9729),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l2101 (
	   .Q (net_6358),
	   .D (n9724),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l2100 (
	   .Q (_net_6174),
	   .D (n9719),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l2099 (
	   .Q (_net_6143),
	   .D (n9714),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l2098 (
	   .Q (_net_6051),
	   .D (n9709),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l2097 (
	   .Q (net_6634),
	   .D (n9704),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l2096 (
	   .Q (_net_5964),
	   .D (n9700),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l2095 (
	   .Q (net_366),
	   .D (n9695),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2094 (
	   .Q (net_6703),
	   .D (n9692),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l2093 (
	   .Q (net_317),
	   .D (n9687),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l2092 (
	   .Q (_net_7560),
	   .D (n9683),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l2091 (
	   .Q (_net_225),
	   .D (n9678),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l2090 (
	   .Q (_net_7588),
	   .D (n9673),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2089 (
	   .Q (net_368),
	   .D (n9668),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2088 (
	   .Q (_net_7656),
	   .D (n9664),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l2087 (
	   .Q (net_7005),
	   .D (n9660),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l2086 (
	   .Q (_net_7327),
	   .D (n9655),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2085 (
	   .Q (net_7548),
	   .D (n9651),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l2084 (
	   .Q (net_7386),
	   .D (n9647),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l2083 (
	   .Q (net_6644),
	   .D (n9642),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l2082 (
	   .Q (_net_7414),
	   .D (n9638),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l2081 (
	   .Q (_net_7436),
	   .D (n9633),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l2080 (
	   .Q (_net_6219),
	   .D (n9628),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l2079 (
	   .Q (net_7205),
	   .D (n9624),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l2078 (
	   .Q (net_6785),
	   .D (n9620),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2077 (
	   .Q (_net_6052),
	   .D (n9616),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l2076 (
	   .Q (net_6307),
	   .D (n9611),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l2075 (
	   .Q (net_6818),
	   .D (n9606),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2074 (
	   .Q (_net_7324),
	   .D (n9602),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2073 (
	   .Q (_net_6153),
	   .D (n9597),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l2072 (
	   .Q (net_6036),
	   .D (n9592),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l2071 (
	   .Q (net_6455),
	   .D (n9588),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l2070 (
	   .Q (_net_7506),
	   .D (n9583),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l2069 (
	   .Q (net_6840),
	   .D (n9579),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l2068 (
	   .Q (net_297),
	   .D (n9574),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l2067 (
	   .Q (_net_7509),
	   .D (n9569),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l2066 (
	   .Q (_net_6021),
	   .D (n9564),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l2065 (
	   .Q (_net_190),
	   .D (n9559),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l2064 (
	   .Q (net_6058),
	   .D (n9554),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l2063 (
	   .Q (net_7524),
	   .D (n9549),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l2062 (
	   .Q (x138),
	   .D (n9546),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l2061 (
	   .Q (net_7183),
	   .D (n9541),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l2060 (
	   .Q (net_6782),
	   .D (n9537),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2059 (
	   .Q (_net_217),
	   .D (n9533),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l2058 (
	   .Q (net_6667),
	   .D (n9528),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l2057 (
	   .Q (net_7015),
	   .D (n9525),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2056 (
	   .Q (net_316),
	   .D (n9520),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l2055 (
	   .Q (net_6871),
	   .D (n9517),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2054 (
	   .Q (_net_7616),
	   .D (n9512),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2053 (
	   .Q (_net_7617),
	   .D (n9507),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2052 (
	   .Q (net_6359),
	   .D (n9502),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l2051 (
	   .Q (_net_7597),
	   .D (n9497),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2050 (
	   .Q (_net_7282),
	   .D (n9492),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2049 (
	   .Q (_net_7415),
	   .D (n9487),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l2048 (
	   .Q (net_6611),
	   .D (n9483),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l2047 (
	   .Q (net_7464),
	   .D (n9478),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l2046 (
	   .Q (net_6842),
	   .D (n9475),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2045 (
	   .Q (net_359),
	   .D (n9470),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l2044 (
	   .Q (net_6972),
	   .D (n9467),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l2043 (
	   .Q (net_6916),
	   .D (n9462),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l2042 (
	   .Q (net_7709),
	   .D (n9459),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l2041 (
	   .Q (_net_6005),
	   .D (n9454),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l2040 (
	   .Q (_net_6280),
	   .D (n9449),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l2039 (
	   .Q (net_6731),
	   .D (n9445),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l2038 (
	   .Q (x638),
	   .D (n9441),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l2037 (
	   .Q (_net_7745),
	   .D (n9436),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l2036 (
	   .Q (net_6775),
	   .D (n9431),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l2035 (
	   .Q (net_145),
	   .D (n9428),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l2034 (
	   .Q (net_6459),
	   .D (n9425),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l2033 (
	   .Q (_net_7317),
	   .D (n9420),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2032 (
	   .Q (_net_6085),
	   .D (n9415),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l2031 (
	   .Q (_net_7569),
	   .D (n9410),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l2030 (
	   .Q (net_6908),
	   .D (n9405),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l2029 (
	   .Q (x0),
	   .D (n9402),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l2028 (
	   .Q (net_6278),
	   .D (n9398),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l2027 (
	   .Q (net_6936),
	   .D (n9393),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l2026 (
	   .Q (net_6601),
	   .D (n9390),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l2025 (
	   .Q (net_7072),
	   .D (n9385),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l2024 (
	   .Q (net_6921),
	   .D (n9381),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2023 (
	   .Q (net_6817),
	   .D (n9377),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2022 (
	   .Q (net_6640),
	   .D (n9373),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2021 (
	   .Q (net_7099),
	   .D (n9370),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l2020 (
	   .Q (net_6265),
	   .D (n9365),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l2019 (
	   .Q (net_6464),
	   .D (n9361),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l2018 (
	   .Q (net_7164),
	   .D (n9356),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l2017 (
	   .Q (_net_7504),
	   .D (n9352),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l2016 (
	   .Q (net_7541),
	   .D (n9348),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l2015 (
	   .Q (net_6535),
	   .D (n9343),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2014 (
	   .Q (net_6662),
	   .D (n9339),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l2013 (
	   .Q (_net_7725),
	   .D (n9335),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l2012 (
	   .Q (_net_5983),
	   .D (n9330),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2011 (
	   .Q (net_6749),
	   .D (n9326),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l2010 (
	   .Q (net_219),
	   .D (n9321),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l2009 (
	   .Q (net_7377),
	   .D (n9316),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l2008 (
	   .Q (_net_7726),
	   .D (n9312),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l2007 (
	   .Q (_net_7516),
	   .D (n9307),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l2006 (
	   .Q (net_7519),
	   .D (n9302),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l2005 (
	   .Q (net_7612),
	   .D (n9298),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2004 (
	   .Q (net_7218),
	   .D (n9294),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l2003 (
	   .Q (net_7190),
	   .D (n9290),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l2002 (
	   .Q (net_6848),
	   .D (n9287),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l2001 (
	   .Q (_net_6137),
	   .D (n9282),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l2000 (
	   .Q (_net_6106),
	   .D (n9277),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1999 (
	   .Q (_net_7530),
	   .D (n9272),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1998 (
	   .Q (net_6669),
	   .D (n9267),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1997 (
	   .Q (_net_7515),
	   .D (n9263),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1996 (
	   .Q (_net_6405),
	   .D (n9258),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1995 (
	   .Q (net_7103),
	   .D (n9254),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1994 (
	   .Q (net_6701),
	   .D (n9250),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1993 (
	   .Q (net_6527),
	   .D (n9245),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1992 (
	   .Q (net_6483),
	   .D (n9242),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1991 (
	   .Q (net_6705),
	   .D (n9238),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1990 (
	   .Q (_net_7701),
	   .D (n9233),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1989 (
	   .Q (net_7463),
	   .D (n9228),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1988 (
	   .Q (net_7156),
	   .D (n9225),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1987 (
	   .Q (_net_6094),
	   .D (n9220),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1986 (
	   .Q (net_7367),
	   .D (n9215),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1985 (
	   .Q (net_7776),
	   .D (n9211),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1984 (
	   .Q (_net_5986),
	   .D (n9206),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1983 (
	   .Q (_net_7682),
	   .D (n9201),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1982 (
	   .Q (net_328),
	   .D (n9196),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1981 (
	   .Q (_net_172),
	   .D (n9192),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1980 (
	   .Q (_net_7260),
	   .D (n9187),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1979 (
	   .Q (net_6492),
	   .D (n9182),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1978 (
	   .Q (net_6253),
	   .D (n9178),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1977 (
	   .Q (_net_6188),
	   .D (n9173),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1976 (
	   .Q (net_6565),
	   .D (n9169),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1975 (
	   .Q (net_6911),
	   .D (n9164),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1974 (
	   .Q (net_318),
	   .D (n9160),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1973 (
	   .Q (_net_7259),
	   .D (n9156),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1972 (
	   .Q (net_162),
	   .D (n9151),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1971 (
	   .Q (net_6665),
	   .D (n9146),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1970 (
	   .Q (net_6876),
	   .D (n9143),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1969 (
	   .Q (net_6520),
	   .D (n9138),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1968 (
	   .Q (net_6333),
	   .D (n9134),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1967 (
	   .Q (_net_7660),
	   .D (n9129),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1966 (
	   .Q (_net_7558),
	   .D (n9124),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1965 (
	   .Q (net_7155),
	   .D (n9120),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1964 (
	   .Q (_net_292),
	   .D (n9115),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1963 (
	   .Q (_net_7804),
	   .D (n9110),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1962 (
	   .Q (_net_7716),
	   .D (n9106),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1961 (
	   .Q (_net_289),
	   .D (n9101),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1960 (
	   .Q (net_256),
	   .D (n9096),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1959 (
	   .Q (net_6270),
	   .D (n9091),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1958 (
	   .Q (net_6649),
	   .D (n9086),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1957 (
	   .Q (net_7084),
	   .D (n9082),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1956 (
	   .Q (net_7101),
	   .D (n9079),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1955 (
	   .Q (_net_115),
	   .D (n9074),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1954 (
	   .Q (net_6306),
	   .D (n9069),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1953 (
	   .Q (net_6984),
	   .D (n9065),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1952 (
	   .Q (net_7305),
	   .D (n9060),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1951 (
	   .Q (net_6966),
	   .D (n9057),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1950 (
	   .Q (_net_7423),
	   .D (n9052),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1949 (
	   .Q (net_7762),
	   .D (n9047),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1948 (
	   .Q (net_230),
	   .D (n9042),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1947 (
	   .Q (net_6937),
	   .D (n9037),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1946 (
	   .Q (net_6864),
	   .D (n9034),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1945 (
	   .Q (x249),
	   .D (n9030),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1944 (
	   .Q (net_6932),
	   .D (n9025),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1943 (
	   .Q (net_6445),
	   .D (n9022),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1942 (
	   .Q (net_6230),
	   .D (n9017),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1941 (
	   .Q (net_7017),
	   .D (n9014),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1940 (
	   .Q (net_6582),
	   .D (n9010),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1939 (
	   .Q (_net_7783),
	   .D (n9005),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1938 (
	   .Q (_net_268),
	   .D (n9000),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1937 (
	   .Q (_net_293),
	   .D (n8995),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1936 (
	   .Q (net_304),
	   .D (n8990),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1935 (
	   .Q (_net_7581),
	   .D (n8986),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1934 (
	   .Q (net_6350),
	   .D (n8981),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1933 (
	   .Q (_net_7466),
	   .D (n8976),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1932 (
	   .Q (net_6534),
	   .D (n8971),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1931 (
	   .Q (_net_209),
	   .D (n8967),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1930 (
	   .Q (net_7544),
	   .D (n8963),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1929 (
	   .Q (net_6326),
	   .D (n8958),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1928 (
	   .Q (_net_7451),
	   .D (n8953),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1927 (
	   .Q (_net_7322),
	   .D (n8948),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1926 (
	   .Q (net_6262),
	   .D (n8943),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1925 (
	   .Q (net_6458),
	   .D (n8939),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1924 (
	   .Q (net_7368),
	   .D (n8934),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1923 (
	   .Q (net_7243),
	   .D (n8931),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1922 (
	   .Q (net_6504),
	   .D (n8926),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1921 (
	   .Q (_net_7787),
	   .D (n8922),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1920 (
	   .Q (_net_6166),
	   .D (n8917),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1919 (
	   .Q (net_6531),
	   .D (n8912),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1918 (
	   .Q (net_6315),
	   .D (n8908),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1917 (
	   .Q (net_6549),
	   .D (n8903),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1916 (
	   .Q (net_7302),
	   .D (n8899),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1915 (
	   .Q (_net_6298),
	   .D (n8895),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1914 (
	   .Q (net_7132),
	   .D (n8891),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1913 (
	   .Q (net_7086),
	   .D (n8886),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1912 (
	   .Q (net_6196),
	   .D (n8882),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1911 (
	   .Q (net_307),
	   .D (n8877),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1910 (
	   .Q (net_6217),
	   .D (n8873),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1909 (
	   .Q (_net_6186),
	   .D (n8869),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1908 (
	   .Q (_net_7806),
	   .D (n8864),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1907 (
	   .Q (_net_7625),
	   .D (n8860),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1906 (
	   .Q (_net_7363),
	   .D (n8855),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1905 (
	   .Q (_net_228),
	   .D (n8850),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1904 (
	   .Q (_net_6048),
	   .D (n8845),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1903 (
	   .Q (_net_7664),
	   .D (n8840),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1902 (
	   .Q (net_7046),
	   .D (n8835),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1901 (
	   .Q (net_195),
	   .D (n8831),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1900 (
	   .Q (net_6787),
	   .D (n8826),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1899 (
	   .Q (net_7542),
	   .D (n8823),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1898 (
	   .Q (_net_7409),
	   .D (n8818),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1897 (
	   .Q (net_7064),
	   .D (n8813),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1896 (
	   .Q (net_6417),
	   .D (n8809),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1895 (
	   .Q (net_6982),
	   .D (n8805),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1894 (
	   .Q (net_7043),
	   .D (n8800),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1893 (
	   .Q (net_6457),
	   .D (n8797),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1892 (
	   .Q (net_6882),
	   .D (n8793),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1891 (
	   .Q (net_6046),
	   .D (n8788),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1890 (
	   .Q (_net_7818),
	   .D (n8784),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1889 (
	   .Q (_net_7265),
	   .D (n8780),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1888 (
	   .Q (_net_7230),
	   .D (n8775),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1887 (
	   .Q (net_387),
	   .D (n8771),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1886 (
	   .Q (net_7110),
	   .D (n8767),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1885 (
	   .Q (_net_6289),
	   .D (n8762),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1884 (
	   .Q (net_6234),
	   .D (n8757),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1883 (
	   .Q (_net_7585),
	   .D (n8753),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1882 (
	   .Q (_net_7476),
	   .D (n8748),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1881 (
	   .Q (_net_6043),
	   .D (n8743),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1880 (
	   .Q (net_7389),
	   .D (n8739),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1879 (
	   .Q (net_7340),
	   .D (n8734),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1878 (
	   .Q (_net_6109),
	   .D (n8730),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1877 (
	   .Q (_net_6824),
	   .D (n8725),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1876 (
	   .Q (_net_7477),
	   .D (n8720),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1875 (
	   .Q (net_333),
	   .D (n8715),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1874 (
	   .Q (net_7521),
	   .D (n8711),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1873 (
	   .Q (x538),
	   .D (n8708),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1872 (
	   .Q (_net_6010),
	   .D (n8703),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1871 (
	   .Q (_net_7811),
	   .D (n8698),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1870 (
	   .Q (_net_6144),
	   .D (n8694),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1869 (
	   .Q (_net_7627),
	   .D (n8689),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1868 (
	   .Q (net_6722),
	   .D (n8685),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1867 (
	   .Q (net_6891),
	   .D (n8681),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1866 (
	   .Q (_net_6418),
	   .D (n8676),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1865 (
	   .Q (_net_7267),
	   .D (n8671),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1864 (
	   .Q (net_7373),
	   .D (n8666),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1863 (
	   .Q (net_198),
	   .D (n8662),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1862 (
	   .Q (net_6600),
	   .D (n8658),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1861 (
	   .Q (net_6577),
	   .D (n8654),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1860 (
	   .Q (net_6865),
	   .D (n8650),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1859 (
	   .Q (_net_6141),
	   .D (n8645),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1858 (
	   .Q (net_6756),
	   .D (n8641),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1857 (
	   .Q (net_6013),
	   .D (n8637),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1856 (
	   .Q (net_6683),
	   .D (n8632),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1855 (
	   .Q (net_151),
	   .D (n8628),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1854 (
	   .Q (net_388),
	   .D (n8625),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1853 (
	   .Q (net_6831),
	   .D (n8621),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1852 (
	   .Q (net_6360),
	   .D (n8616),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1851 (
	   .Q (net_6463),
	   .D (n8612),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1850 (
	   .Q (net_181),
	   .D (n8607),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1849 (
	   .Q (_net_7319),
	   .D (n8602),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1848 (
	   .Q (net_6695),
	   .D (n8598),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1847 (
	   .Q (_net_7695),
	   .D (n8593),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1846 (
	   .Q (net_7778),
	   .D (n8588),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1845 (
	   .Q (_net_6282),
	   .D (n8583),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1844 (
	   .Q (net_350),
	   .D (n8578),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1843 (
	   .Q (net_6475),
	   .D (n8575),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1842 (
	   .Q (_net_122),
	   .D (n8570),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1841 (
	   .Q (net_6794),
	   .D (n8565),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1840 (
	   .Q (net_6956),
	   .D (n8561),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1839 (
	   .Q (net_166),
	   .D (n8557),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1838 (
	   .Q (net_6792),
	   .D (n8552),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1837 (
	   .Q (net_6707),
	   .D (n8549),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1836 (
	   .Q (net_6499),
	   .D (n8544),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1835 (
	   .Q (net_239),
	   .D (n8540),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1834 (
	   .Q (net_6771),
	   .D (n8535),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1833 (
	   .Q (_net_7284),
	   .D (n8531),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1832 (
	   .Q (_net_7349),
	   .D (n8526),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1831 (
	   .Q (net_6838),
	   .D (n8522),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1830 (
	   .Q (_net_7575),
	   .D (n8517),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1829 (
	   .Q (net_6744),
	   .D (n8513),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1828 (
	   .Q (_net_6557),
	   .D (n8508),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1827 (
	   .Q (net_6622),
	   .D (n8504),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1826 (
	   .Q (_net_6039),
	   .D (n8499),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1825 (
	   .Q (net_7212),
	   .D (n8494),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1824 (
	   .Q (net_7020),
	   .D (n8491),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1823 (
	   .Q (_net_6178),
	   .D (n8486),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1822 (
	   .Q (_net_7450),
	   .D (n8481),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1821 (
	   .Q (net_6754),
	   .D (n8477),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1820 (
	   .Q (_net_5961),
	   .D (n8472),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1819 (
	   .Q (net_7039),
	   .D (n8467),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1818 (
	   .Q (net_6742),
	   .D (n8464),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1817 (
	   .Q (net_6518),
	   .D (n8459),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1816 (
	   .Q (net_6945),
	   .D (n8455),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1815 (
	   .Q (net_7459),
	   .D (n8451),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1814 (
	   .Q (net_7375),
	   .D (n8447),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1813 (
	   .Q (_net_7687),
	   .D (n8443),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1812 (
	   .Q (_net_5924),
	   .D (n8438),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1811 (
	   .Q (x342),
	   .D (n8435),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1810 (
	   .Q (net_332),
	   .D (n8430),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1809 (
	   .Q (_net_6089),
	   .D (n8426),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1808 (
	   .Q (net_7237),
	   .D (n8422),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1807 (
	   .Q (net_6393),
	   .D (n8418),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1806 (
	   .Q (net_7137),
	   .D (n8415),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1805 (
	   .Q (_net_7333),
	   .D (n8410),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1804 (
	   .Q (_net_6958),
	   .D (n8405),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1803 (
	   .Q (net_7104),
	   .D (n8401),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1802 (
	   .Q (_net_7568),
	   .D (n8396),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1801 (
	   .Q (net_6425),
	   .D (n8392),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1800 (
	   .Q (_net_6027),
	   .D (n8387),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1799 (
	   .Q (_net_7602),
	   .D (n8382),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1798 (
	   .Q (_net_7735),
	   .D (n8377),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1797 (
	   .Q (_net_7685),
	   .D (n8372),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1796 (
	   .Q (_net_189),
	   .D (n8367),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1795 (
	   .Q (net_7605),
	   .D (n8362),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1794 (
	   .Q (net_6427),
	   .D (n8359),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1793 (
	   .Q (_net_6823),
	   .D (n8354),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1792 (
	   .Q (net_7023),
	   .D (n8350),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1791 (
	   .Q (_net_6123),
	   .D (n8345),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1790 (
	   .Q (net_6809),
	   .D (n8340),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1789 (
	   .Q (net_143),
	   .D (n8337),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1788 (
	   .Q (net_6851),
	   .D (n8334),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1787 (
	   .Q (net_6276),
	   .D (n8329),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1786 (
	   .Q (_net_6201),
	   .D (n8324),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1785 (
	   .Q (net_7138),
	   .D (n8320),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1784 (
	   .Q (net_6853),
	   .D (n8316),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1783 (
	   .Q (net_7186),
	   .D (n8311),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1782 (
	   .Q (net_7181),
	   .D (n8307),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1781 (
	   .Q (net_7045),
	   .D (n8303),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1780 (
	   .Q (_net_6020),
	   .D (n8299),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1779 (
	   .Q (_net_7648),
	   .D (n8294),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1778 (
	   .Q (net_6321),
	   .D (n8289),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1777 (
	   .Q (_net_6413),
	   .D (n8284),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1776 (
	   .Q (net_7538),
	   .D (n8280),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1775 (
	   .Q (net_6615),
	   .D (n8276),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1774 (
	   .Q (net_6312),
	   .D (n8271),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1773 (
	   .Q (net_7169),
	   .D (n8266),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1772 (
	   .Q (net_7615),
	   .D (n8262),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1771 (
	   .Q (net_196),
	   .D (n8258),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1770 (
	   .Q (_net_7432),
	   .D (n8253),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1769 (
	   .Q (net_6389),
	   .D (n8249),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1768 (
	   .Q (net_6494),
	   .D (n8245),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1767 (
	   .Q (net_370),
	   .D (n8241),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1766 (
	   .Q (_net_7580),
	   .D (n8237),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1765 (
	   .Q (net_7177),
	   .D (n8232),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1764 (
	   .Q (net_6910),
	   .D (n8228),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1763 (
	   .Q (_net_7755),
	   .D (n8224),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1762 (
	   .Q (net_6390),
	   .D (n8220),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1761 (
	   .Q (_net_7702),
	   .D (n8216),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1760 (
	   .Q (net_7772),
	   .D (n8211),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1759 (
	   .Q (net_6678),
	   .D (n8206),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1758 (
	   .Q (_net_6159),
	   .D (n8202),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1757 (
	   .Q (net_275),
	   .D (n8197),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1756 (
	   .Q (_net_7275),
	   .D (n8192),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1755 (
	   .Q (net_6835),
	   .D (n8188),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1754 (
	   .Q (net_6767),
	   .D (n8183),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1753 (
	   .Q (_net_180),
	   .D (n8179),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1752 (
	   .Q (net_6682),
	   .D (n8174),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1751 (
	   .Q (_net_221),
	   .D (n8170),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1750 (
	   .Q (net_7715),
	   .D (n8166),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1749 (
	   .Q (net_242),
	   .D (n8161),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1748 (
	   .Q (net_7339),
	   .D (n8156),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1747 (
	   .Q (_net_262),
	   .D (n8152),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1746 (
	   .Q (net_6638),
	   .D (n8147),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1745 (
	   .Q (net_6571),
	   .D (n8144),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1744 (
	   .Q (net_7141),
	   .D (n8140),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1743 (
	   .Q (_net_7592),
	   .D (n8135),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1742 (
	   .Q (_net_7291),
	   .D (n8130),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1741 (
	   .Q (net_6895),
	   .D (n8125),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1740 (
	   .Q (_net_7562),
	   .D (n8121),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1739 (
	   .Q (net_6798),
	   .D (n8116),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1738 (
	   .Q (_net_6115),
	   .D (n8112),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1737 (
	   .Q (_net_7417),
	   .D (n8107),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1736 (
	   .Q (_net_7499),
	   .D (n8102),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1735 (
	   .Q (_net_7573),
	   .D (n8097),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1734 (
	   .Q (net_7036),
	   .D (n8092),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1733 (
	   .Q (net_285),
	   .D (n8088),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1732 (
	   .Q (net_6596),
	   .D (n8085),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1731 (
	   .Q (_net_7262),
	   .D (n8080),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1730 (
	   .Q (net_6924),
	   .D (n8075),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1729 (
	   .Q (net_6614),
	   .D (n8072),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1728 (
	   .Q (net_6675),
	   .D (n8067),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1727 (
	   .Q (net_6968),
	   .D (n8064),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1726 (
	   .Q (net_6919),
	   .D (n8059),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1725 (
	   .Q (net_6988),
	   .D (n8056),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1724 (
	   .Q (net_344),
	   .D (n8051),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1723 (
	   .Q (net_6365),
	   .D (n8047),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1722 (
	   .Q (net_7744),
	   .D (n8042),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1721 (
	   .Q (net_7680),
	   .D (n8038),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1720 (
	   .Q (_net_6072),
	   .D (n8033),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1719 (
	   .Q (net_6542),
	   .D (n8028),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1718 (
	   .Q (_net_6287),
	   .D (n8024),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1717 (
	   .Q (_net_291),
	   .D (n8019),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1716 (
	   .Q (net_7131),
	   .D (n8015),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1715 (
	   .Q (_net_5852),
	   .D (n8010),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1714 (
	   .Q (net_379),
	   .D (n8005),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1713 (
	   .Q (net_6975),
	   .D (n8002),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1712 (
	   .Q (net_7087),
	   .D (n7997),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1711 (
	   .Q (net_6585),
	   .D (n7994),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1710 (
	   .Q (net_6651),
	   .D (n7989),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1709 (
	   .Q (_net_7425),
	   .D (n7985),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1708 (
	   .Q (net_158),
	   .D (n7980),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1707 (
	   .Q (_net_5855),
	   .D (n7975),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1706 (
	   .Q (net_7491),
	   .D (n7970),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1705 (
	   .Q (net_6992),
	   .D (n7967),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1704 (
	   .Q (net_7078),
	   .D (n7962),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1703 (
	   .Q (net_6232),
	   .D (n7958),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1702 (
	   .Q (net_6724),
	   .D (n7955),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1701 (
	   .Q (net_6056),
	   .D (n7950),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1700 (
	   .Q (net_335),
	   .D (n7945),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1699 (
	   .Q (net_7540),
	   .D (n7942),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1698 (
	   .Q (net_6930),
	   .D (n7937),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1697 (
	   .Q (net_237),
	   .D (n7933),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1696 (
	   .Q (net_6568),
	   .D (n7929),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1695 (
	   .Q (net_7456),
	   .D (n7924),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1694 (
	   .Q (net_311),
	   .D (n7920),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1693 (
	   .Q (net_6363),
	   .D (n7916),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1692 (
	   .Q (_net_6552),
	   .D (n7911),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1691 (
	   .Q (net_7192),
	   .D (n7906),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1690 (
	   .Q (_net_6031),
	   .D (n7902),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1689 (
	   .Q (_net_5850),
	   .D (n7897),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1688 (
	   .Q (net_7249),
	   .D (n7893),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1687 (
	   .Q (_net_7484),
	   .D (n7888),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1686 (
	   .Q (net_6344),
	   .D (n7883),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1685 (
	   .Q (net_7673),
	   .D (n7878),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1684 (
	   .Q (net_6874),
	   .D (n7875),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1683 (
	   .Q (net_137),
	   .D (n7871),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1682 (
	   .Q (net_358),
	   .D (n7867),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1681 (
	   .Q (_net_6409),
	   .D (n7863),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1680 (
	   .Q (_net_5971),
	   .D (n7858),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1679 (
	   .Q (net_200),
	   .D (n7853),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1678 (
	   .Q (net_327),
	   .D (n7848),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1677 (
	   .Q (x264),
	   .D (n7845),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1676 (
	   .Q (net_6331),
	   .D (n7840),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1675 (
	   .Q (_net_7276),
	   .D (n7835),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1674 (
	   .Q (net_6566),
	   .D (n7831),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1673 (
	   .Q (net_6528),
	   .D (n7826),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1672 (
	   .Q (_net_5974),
	   .D (n7822),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1671 (
	   .Q (net_6387),
	   .D (n7818),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1670 (
	   .Q (net_6734),
	   .D (n7815),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1669 (
	   .Q (net_6659),
	   .D (n7810),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1668 (
	   .Q (net_6947),
	   .D (n7806),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1667 (
	   .Q (net_6797),
	   .D (n7802),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1666 (
	   .Q (_net_7442),
	   .D (n7798),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1665 (
	   .Q (_net_6049),
	   .D (n7793),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1664 (
	   .Q (_net_6093),
	   .D (n7788),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1663 (
	   .Q (net_6710),
	   .D (n7784),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1662 (
	   .Q (net_7059),
	   .D (n7779),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1661 (
	   .Q (net_6397),
	   .D (n7776),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1660 (
	   .Q (x420),
	   .D (n7773),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1659 (
	   .Q (_net_7699),
	   .D (n7768),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1658 (
	   .Q (net_7160),
	   .D (n7764),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1657 (
	   .Q (net_7143),
	   .D (n7760),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1656 (
	   .Q (net_6441),
	   .D (n7756),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1655 (
	   .Q (_net_7555),
	   .D (n7751),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1654 (
	   .Q (_net_6828),
	   .D (n7746),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1653 (
	   .Q (_net_392),
	   .D (n7741),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1652 (
	   .Q (x522),
	   .D (n7737),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1651 (
	   .Q (net_7526),
	   .D (n7732),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1650 (
	   .Q (_net_7289),
	   .D (n7728),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1649 (
	   .Q (_net_7273),
	   .D (n7723),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1648 (
	   .Q (net_6837),
	   .D (n7719),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1647 (
	   .Q (net_7764),
	   .D (n7714),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1646 (
	   .Q (net_6047),
	   .D (n7709),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1645 (
	   .Q (net_6304),
	   .D (n7704),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1644 (
	   .Q (net_6748),
	   .D (n7700),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1643 (
	   .Q (_net_5995),
	   .D (n7695),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1642 (
	   .Q (x38),
	   .D (n7691),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1641 (
	   .Q (net_231),
	   .D (n7686),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1640 (
	   .Q (_net_125),
	   .D (n7681),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1639 (
	   .Q (_net_6103),
	   .D (n7676),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1638 (
	   .Q (_net_6091),
	   .D (n7671),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1637 (
	   .Q (_net_7228),
	   .D (n7666),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1636 (
	   .Q (net_7486),
	   .D (n7661),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1635 (
	   .Q (net_6467),
	   .D (n7658),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1634 (
	   .Q (net_7139),
	   .D (n7654),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1633 (
	   .Q (net_6299),
	   .D (n7649),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1632 (
	   .Q (net_341),
	   .D (n7644),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1631 (
	   .Q (_net_5999),
	   .D (n7640),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1630 (
	   .Q (net_7668),
	   .D (n7635),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1629 (
	   .Q (_net_7331),
	   .D (n7631),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1628 (
	   .Q (net_7489),
	   .D (n7626),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1627 (
	   .Q (_net_6207),
	   .D (n7622),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1626 (
	   .Q (net_7392),
	   .D (n7618),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1625 (
	   .Q (net_199),
	   .D (n7613),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1624 (
	   .Q (_net_6959),
	   .D (n7608),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1623 (
	   .Q (net_6716),
	   .D (n7604),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1622 (
	   .Q (net_7494),
	   .D (n7599),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1621 (
	   .Q (x187),
	   .D (n7596),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1620 (
	   .Q (_net_127),
	   .D (n7591),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1619 (
	   .Q (_net_6033),
	   .D (n7586),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1618 (
	   .Q (net_6811),
	   .D (n7581),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1617 (
	   .Q (_net_6319),
	   .D (n7577),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1616 (
	   .Q (_net_6127),
	   .D (n7572),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1615 (
	   .Q (_net_7824),
	   .D (n7567),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1614 (
	   .Q (_net_7293),
	   .D (n7563),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1613 (
	   .Q (_net_7381),
	   .D (n7558),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1612 (
	   .Q (net_6266),
	   .D (n7553),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1611 (
	   .Q (net_243),
	   .D (n7548),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1610 (
	   .Q (_net_177),
	   .D (n7543),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1609 (
	   .Q (x476),
	   .D (n7539),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1608 (
	   .Q (net_6757),
	   .D (n7535),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1607 (
	   .Q (net_7210),
	   .D (n7530),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1606 (
	   .Q (net_6451),
	   .D (n7527),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1605 (
	   .Q (net_7211),
	   .D (n7522),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1604 (
	   .Q (_net_7471),
	   .D (n7518),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1603 (
	   .Q (net_6550),
	   .D (n7513),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1602 (
	   .Q (net_6774),
	   .D (n7509),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1601 (
	   .Q (net_348),
	   .D (n7505),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1600 (
	   .Q (_net_264),
	   .D (n7501),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1599 (
	   .Q (_net_6068),
	   .D (n7496),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1598 (
	   .Q (net_6726),
	   .D (n7492),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1597 (
	   .Q (_net_6962),
	   .D (n7487),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1596 (
	   .Q (net_7077),
	   .D (n7482),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1595 (
	   .Q (_net_7351),
	   .D (n7478),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1594 (
	   .Q (_net_6222),
	   .D (n7473),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1593 (
	   .Q (net_6337),
	   .D (n7468),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1592 (
	   .Q (net_7216),
	   .D (n7463),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1591 (
	   .Q (_net_7263),
	   .D (n7459),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1590 (
	   .Q (_net_6007),
	   .D (n7454),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1589 (
	   .Q (net_6740),
	   .D (n7450),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1588 (
	   .Q (net_6696),
	   .D (n7446),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1587 (
	   .Q (net_6700),
	   .D (n7442),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1586 (
	   .Q (_net_6069),
	   .D (n7437),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1585 (
	   .Q (_net_7757),
	   .D (n7432),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1584 (
	   .Q (net_6345),
	   .D (n7427),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1583 (
	   .Q (_net_6957),
	   .D (n7422),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1582 (
	   .Q (net_6257),
	   .D (n7417),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1581 (
	   .Q (net_6994),
	   .D (n7413),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1580 (
	   .Q (net_7054),
	   .D (n7408),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1579 (
	   .Q (net_6503),
	   .D (n7404),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1578 (
	   .Q (_net_7473),
	   .D (n7400),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1577 (
	   .Q (_net_117),
	   .D (n7395),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1576 (
	   .Q (net_7118),
	   .D (n7391),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1575 (
	   .Q (_net_6105),
	   .D (n7386),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1574 (
	   .Q (_net_7666),
	   .D (n7381),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1573 (
	   .Q (net_6228),
	   .D (n7376),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1572 (
	   .Q (net_7065),
	   .D (n7372),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1571 (
	   .Q (net_6317),
	   .D (n7368),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1570 (
	   .Q (net_185),
	   .D (n7363),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1569 (
	   .Q (net_7008),
	   .D (n7359),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1568 (
	   .Q (net_250),
	   .D (n7354),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1567 (
	   .Q (net_6193),
	   .D (n7349),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1566 (
	   .Q (net_7173),
	   .D (n7344),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1565 (
	   .Q (_net_6179),
	   .D (n7340),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1564 (
	   .Q (net_5860),
	   .D (n7335),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1563 (
	   .Q (net_6264),
	   .D (n7330),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1562 (
	   .Q (net_6715),
	   .D (n7326),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1561 (
	   .Q (_net_7365),
	   .D (n7321),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1560 (
	   .Q (net_6374),
	   .D (n7316),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1559 (
	   .Q (net_6869),
	   .D (n7312),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1558 (
	   .Q (_net_7697),
	   .D (n7307),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1557 (
	   .Q (_net_6288),
	   .D (n7302),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1556 (
	   .Q (_net_6028),
	   .D (n7297),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1555 (
	   .Q (_net_7816),
	   .D (n7292),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1554 (
	   .Q (net_342),
	   .D (n7288),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1553 (
	   .Q (net_6511),
	   .D (n7284),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1552 (
	   .Q (_net_6026),
	   .D (n7280),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1551 (
	   .Q (_net_6291),
	   .D (n7275),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1550 (
	   .Q (_net_6151),
	   .D (n7270),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1549 (
	   .Q (_net_6402),
	   .D (n7265),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1548 (
	   .Q (net_6627),
	   .D (n7260),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1547 (
	   .Q (_net_7791),
	   .D (n7256),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1546 (
	   .Q (net_6801),
	   .D (n7252),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1545 (
	   .Q (net_7807),
	   .D (n7249),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1544 (
	   .Q (_net_6423),
	   .D (n7245),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1543 (
	   .Q (_net_6145),
	   .D (n7240),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1542 (
	   .Q (_net_6295),
	   .D (n7235),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1541 (
	   .Q (net_7090),
	   .D (n7230),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1540 (
	   .Q (_net_6200),
	   .D (n7226),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1539 (
	   .Q (net_6211),
	   .D (n7221),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1538 (
	   .Q (_net_7361),
	   .D (n7216),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1537 (
	   .Q (net_6559),
	   .D (n7212),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1536 (
	   .Q (_net_6080),
	   .D (n7207),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1535 (
	   .Q (net_6477),
	   .D (n7203),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1534 (
	   .Q (net_7238),
	   .D (n7199),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1533 (
	   .Q (_net_6554),
	   .D (n7194),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1532 (
	   .Q (net_6430),
	   .D (n7190),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1531 (
	   .Q (net_7307),
	   .D (n7185),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1530 (
	   .Q (net_7543),
	   .D (n7182),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1529 (
	   .Q (net_161),
	   .D (n7177),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1528 (
	   .Q (_net_5979),
	   .D (n7172),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1527 (
	   .Q (net_6235),
	   .D (n7167),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1526 (
	   .Q (x195),
	   .D (n7164),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1525 (
	   .Q (net_6862),
	   .D (n7160),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1524 (
	   .Q (net_7226),
	   .D (n7155),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1523 (
	   .Q (net_6948),
	   .D (n7151),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1522 (
	   .Q (net_6249),
	   .D (n7147),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1521 (
	   .Q (net_7496),
	   .D (n7142),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1520 (
	   .Q (_net_5848),
	   .D (n7138),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1519 (
	   .Q (_net_7705),
	   .D (n7133),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1518 (
	   .Q (net_6660),
	   .D (n7128),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1517 (
	   .Q (net_6561),
	   .D (n7125),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1516 (
	   .Q (net_6498),
	   .D (n7120),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1515 (
	   .Q (net_6329),
	   .D (n7116),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1514 (
	   .Q (net_7088),
	   .D (n7111),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1513 (
	   .Q (net_7769),
	   .D (n7107),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1512 (
	   .Q (_net_193),
	   .D (n7102),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1511 (
	   .Q (net_7152),
	   .D (n7098),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1510 (
	   .Q (net_383),
	   .D (n7093),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1509 (
	   .Q (net_6673),
	   .D (n7089),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1508 (
	   .Q (net_7460),
	   .D (n7085),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1507 (
	   .Q (net_6872),
	   .D (n7082),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1506 (
	   .Q (_net_6285),
	   .D (n7077),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1505 (
	   .Q (_net_7761),
	   .D (n7072),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1504 (
	   .Q (_net_6122),
	   .D (n7067),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1503 (
	   .Q (net_6769),
	   .D (n7062),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1502 (
	   .Q (_net_7268),
	   .D (n7058),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1501 (
	   .Q (_net_7579),
	   .D (n7053),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1500 (
	   .Q (net_6394),
	   .D (n7049),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1499 (
	   .Q (net_6378),
	   .D (n7045),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1498 (
	   .Q (net_6889),
	   .D (n7041),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1497 (
	   .Q (net_306),
	   .D (n7036),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1496 (
	   .Q (_net_7298),
	   .D (n7032),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1495 (
	   .Q (net_6902),
	   .D (n7027),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1494 (
	   .Q (net_222),
	   .D (n7023),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1493 (
	   .Q (_net_6140),
	   .D (n7018),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1492 (
	   .Q (_net_7408),
	   .D (n7013),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1491 (
	   .Q (net_6597),
	   .D (n7009),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1490 (
	   .Q (net_6621),
	   .D (n7005),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1489 (
	   .Q (_net_281),
	   .D (n7000),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1488 (
	   .Q (_net_7256),
	   .D (n6995),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1487 (
	   .Q (net_6495),
	   .D (n6990),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1486 (
	   .Q (net_7172),
	   .D (n6986),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1485 (
	   .Q (net_6342),
	   .D (n6982),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1484 (
	   .Q (net_7051),
	   .D (n6977),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1483 (
	   .Q (net_7245),
	   .D (n6974),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1482 (
	   .Q (net_194),
	   .D (n6969),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1481 (
	   .Q (_net_6098),
	   .D (n6964),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1480 (
	   .Q (net_149),
	   .D (n6960),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1479 (
	   .Q (net_6587),
	   .D (n6957),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1478 (
	   .Q (_net_7500),
	   .D (n6952),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1477 (
	   .Q (net_375),
	   .D (n6947),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1476 (
	   .Q (_net_7589),
	   .D (n6943),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1475 (
	   .Q (_net_114),
	   .D (n6938),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1474 (
	   .Q (net_7150),
	   .D (n6934),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1473 (
	   .Q (net_244),
	   .D (n6929),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1472 (
	   .Q (_net_7443),
	   .D (n6924),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1471 (
	   .Q (net_7309),
	   .D (n6919),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1470 (
	   .Q (_net_215),
	   .D (n6915),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1469 (
	   .Q (net_7053),
	   .D (n6910),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1468 (
	   .Q (net_6904),
	   .D (n6906),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1467 (
	   .Q (net_340),
	   .D (n6902),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1466 (
	   .Q (net_6607),
	   .D (n6899),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1465 (
	   .Q (net_7009),
	   .D (n6895),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1464 (
	   .Q (_net_7427),
	   .D (n6890),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1463 (
	   .Q (net_6712),
	   .D (n6886),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1462 (
	   .Q (_net_6161),
	   .D (n6881),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1461 (
	   .Q (net_7209),
	   .D (n6876),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1460 (
	   .Q (net_216),
	   .D (n6872),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1459 (
	   .Q (net_7193),
	   .D (n6867),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1458 (
	   .Q (net_7166),
	   .D (n6863),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1457 (
	   .Q (net_6470),
	   .D (n6860),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1456 (
	   .Q (_net_5990),
	   .D (n6855),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1455 (
	   .Q (net_240),
	   .D (n6850),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1454 (
	   .Q (_net_7325),
	   .D (n6845),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1453 (
	   .Q (_net_5993),
	   .D (n6840),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1452 (
	   .Q (net_7025),
	   .D (n6836),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1451 (
	   .Q (_net_7584),
	   .D (n6831),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1450 (
	   .Q (net_7044),
	   .D (n6826),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1449 (
	   .Q (net_301),
	   .D (n6822),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1448 (
	   .Q (_net_7700),
	   .D (n6818),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1447 (
	   .Q (net_7033),
	   .D (n6813),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1446 (
	   .Q (net_6526),
	   .D (n6809),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1445 (
	   .Q (net_6990),
	   .D (n6806),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1444 (
	   .Q (_net_7258),
	   .D (n6801),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1443 (
	   .Q (net_6933),
	   .D (n6796),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1442 (
	   .Q (net_7394),
	   .D (n6793),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1441 (
	   .Q (_net_7446),
	   .D (n6788),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1440 (
	   .Q (net_6519),
	   .D (n6783),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1439 (
	   .Q (_net_7723),
	   .D (n6779),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1438 (
	   .Q (_net_6117),
	   .D (n6774),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1437 (
	   .Q (net_6830),
	   .D (n6770),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1436 (
	   .Q (_net_6136),
	   .D (n6765),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1435 (
	   .Q (net_6728),
	   .D (n6761),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1434 (
	   .Q (net_314),
	   .D (n6756),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1433 (
	   .Q (net_6894),
	   .D (n6752),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1432 (
	   .Q (net_147),
	   .D (n6749),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1431 (
	   .Q (net_7549),
	   .D (n6746),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1430 (
	   .Q (_net_7620),
	   .D (n6741),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1429 (
	   .Q (net_136),
	   .D (n6736),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1428 (
	   .Q (net_7180),
	   .D (n6732),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1427 (
	   .Q (_net_6113),
	   .D (n6727),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1426 (
	   .Q (net_7345),
	   .D (n6722),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1425 (
	   .Q (net_6793),
	   .D (n6717),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1424 (
	   .Q (net_6655),
	   .D (n6713),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1423 (
	   .Q (_net_7279),
	   .D (n6709),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1422 (
	   .Q (net_7029),
	   .D (n6704),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1421 (
	   .Q (net_6353),
	   .D (n6700),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1420 (
	   .Q (_net_7623),
	   .D (n6695),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1419 (
	   .Q (x681),
	   .D (n6691),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1418 (
	   .Q (net_6997),
	   .D (n6687),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1417 (
	   .Q (_net_278),
	   .D (n6682),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1416 (
	   .Q (net_6708),
	   .D (n6678),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1415 (
	   .Q (net_6834),
	   .D (n6674),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1414 (
	   .Q (net_315),
	   .D (n6669),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1413 (
	   .Q (_net_6129),
	   .D (n6665),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1412 (
	   .Q (net_6424),
	   .D (n6661),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1411 (
	   .Q (net_7638),
	   .D (n6656),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1410 (
	   .Q (_net_124),
	   .D (n6652),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1409 (
	   .Q (net_7145),
	   .D (n6648),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1408 (
	   .Q (net_6003),
	   .D (n6643),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1407 (
	   .Q (net_7187),
	   .D (n6638),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1406 (
	   .Q (_net_6170),
	   .D (n6634),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1405 (
	   .Q (net_6261),
	   .D (n6629),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1404 (
	   .Q (net_168),
	   .D (n6624),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1403 (
	   .Q (net_7163),
	   .D (n6619),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1402 (
	   .Q (net_6917),
	   .D (n6615),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1401 (
	   .Q (net_6272),
	   .D (n6611),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1400 (
	   .Q (_net_5976),
	   .D (n6606),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1399 (
	   .Q (_net_7448),
	   .D (n6601),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1398 (
	   .Q (_net_6119),
	   .D (n6596),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1397 (
	   .Q (net_157),
	   .D (n6591),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1396 (
	   .Q (net_6814),
	   .D (n6586),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1395 (
	   .Q (net_386),
	   .D (n6583),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1394 (
	   .Q (net_6226),
	   .D (n6578),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1393 (
	   .Q (net_7485),
	   .D (n6574),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1392 (
	   .Q (_net_6146),
	   .D (n6570),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1391 (
	   .Q (net_6382),
	   .D (n6566),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1390 (
	   .Q (net_6846),
	   .D (n6563),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1389 (
	   .Q (_net_7654),
	   .D (n6558),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1388 (
	   .Q (net_6713),
	   .D (n6554),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1387 (
	   .Q (net_7397),
	   .D (n6550),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1386 (
	   .Q (_net_118),
	   .D (n6545),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1385 (
	   .Q (_net_6126),
	   .D (n6540),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1384 (
	   .Q (net_7606),
	   .D (n6535),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1383 (
	   .Q (net_330),
	   .D (n6531),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1382 (
	   .Q (_net_5857),
	   .D (n6527),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1381 (
	   .Q (_net_7805),
	   .D (n6522),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1380 (
	   .Q (net_6866),
	   .D (n6519),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1379 (
	   .Q (net_6836),
	   .D (n6515),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1378 (
	   .Q (net_6604),
	   .D (n6511),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1377 (
	   .Q (net_6563),
	   .D (n6507),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1376 (
	   .Q (net_7074),
	   .D (n6502),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1375 (
	   .Q (net_6355),
	   .D (n6498),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1374 (
	   .Q (net_205),
	   .D (n6493),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1373 (
	   .Q (net_7242),
	   .D (n6489),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1372 (
	   .Q (net_6462),
	   .D (n6485),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1371 (
	   .Q (net_6626),
	   .D (n6480),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1370 (
	   .Q (net_7148),
	   .D (n6477),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1369 (
	   .Q (net_6777),
	   .D (n6472),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1368 (
	   .Q (net_6980),
	   .D (n6469),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1367 (
	   .Q (net_6647),
	   .D (n6464),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1366 (
	   .Q (net_6348),
	   .D (n6460),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1365 (
	   .Q (_net_7257),
	   .D (n6455),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1364 (
	   .Q (_net_6692),
	   .D (n6450),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1363 (
	   .Q (net_6702),
	   .D (n6446),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1362 (
	   .Q (net_7069),
	   .D (n6441),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1361 (
	   .Q (net_7462),
	   .D (n6437),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1360 (
	   .Q (net_156),
	   .D (n6432),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1359 (
	   .Q (net_6826),
	   .D (n6427),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1358 (
	   .Q (net_6383),
	   .D (n6423),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1357 (
	   .Q (net_6625),
	   .D (n6419),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1356 (
	   .Q (net_7208),
	   .D (n6415),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1355 (
	   .Q (_net_7438),
	   .D (n6411),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1354 (
	   .Q (net_6481),
	   .D (n6407),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1353 (
	   .Q (net_6738),
	   .D (n6403),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1352 (
	   .Q (net_6399),
	   .D (n6399),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1351 (
	   .Q (_net_6101),
	   .D (n6395),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1350 (
	   .Q (net_6361),
	   .D (n6390),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1349 (
	   .Q (net_7117),
	   .D (n6386),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1348 (
	   .Q (_net_7661),
	   .D (n6381),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1347 (
	   .Q (net_7341),
	   .D (n6376),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1346 (
	   .Q (_net_7098),
	   .D (n6371),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1345 (
	   .Q (net_6439),
	   .D (n6367),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1344 (
	   .Q (_net_7440),
	   .D (n6362),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1343 (
	   .Q (net_6679),
	   .D (n6357),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1342 (
	   .Q (net_6747),
	   .D (n6354),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1341 (
	   .Q (net_131),
	   .D (n6350),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1340 (
	   .Q (_net_7353),
	   .D (n6346),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1339 (
	   .Q (net_6469),
	   .D (n6342),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1338 (
	   .Q (_net_6074),
	   .D (n6337),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1337 (
	   .Q (net_381),
	   .D (n6332),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1336 (
	   .Q (net_7161),
	   .D (n6329),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1335 (
	   .Q (_net_6001),
	   .D (n6324),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1334 (
	   .Q (_net_5922),
	   .D (n6319),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1333 (
	   .Q (net_7770),
	   .D (n6316),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1332 (
	   .Q (_net_5994),
	   .D (n6311),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1331 (
	   .Q (net_302),
	   .D (n6306),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1330 (
	   .Q (net_7454),
	   .D (n6302),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1329 (
	   .Q (net_7130),
	   .D (n6299),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1328 (
	   .Q (_net_7789),
	   .D (n6294),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1327 (
	   .Q (x718),
	   .D (n6290),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1326 (
	   .Q (net_6212),
	   .D (n6285),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1325 (
	   .Q (_net_174),
	   .D (n6281),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1324 (
	   .Q (net_7752),
	   .D (n6276),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1323 (
	   .Q (net_167),
	   .D (n6271),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1322 (
	   .Q (_net_7434),
	   .D (n6266),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1321 (
	   .Q (_net_7801),
	   .D (n6261),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1320 (
	   .Q (net_6750),
	   .D (n6258),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1319 (
	   .Q (net_6697),
	   .D (n6254),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1318 (
	   .Q (_net_201),
	   .D (n6249),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1317 (
	   .Q (_net_210),
	   .D (n6244),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1316 (
	   .Q (net_385),
	   .D (n6239),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1315 (
	   .Q (net_6629),
	   .D (n6235),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1314 (
	   .Q (net_7739),
	   .D (n6231),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1313 (
	   .Q (net_186),
	   .D (n6227),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1312 (
	   .Q (net_7679),
	   .D (n6222),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1311 (
	   .Q (_net_6099),
	   .D (n6218),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1310 (
	   .Q (net_7385),
	   .D (n6214),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1309 (
	   .Q (_net_7254),
	   .D (n6209),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1308 (
	   .Q (net_382),
	   .D (n6204),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1307 (
	   .Q (_net_7693),
	   .D (n6200),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1306 (
	   .Q (net_6508),
	   .D (n6195),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1305 (
	   .Q (_net_6149),
	   .D (n6191),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1304 (
	   .Q (_net_6124),
	   .D (n6186),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1303 (
	   .Q (net_6309),
	   .D (n6181),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1302 (
	   .Q (net_6301),
	   .D (n6176),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1301 (
	   .Q (_net_6071),
	   .D (n6171),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1300 (
	   .Q (_net_6209),
	   .D (n6166),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1299 (
	   .Q (net_7083),
	   .D (n6161),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1298 (
	   .Q (net_6892),
	   .D (n6158),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1297 (
	   .Q (_net_6293),
	   .D (n6153),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1296 (
	   .Q (net_274),
	   .D (n6148),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1295 (
	   .Q (net_6594),
	   .D (n6145),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1294 (
	   .Q (_net_7681),
	   .D (n6140),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1293 (
	   .Q (net_6385),
	   .D (n6136),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1292 (
	   .Q (_net_7808),
	   .D (n6132),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1291 (
	   .Q (net_7038),
	   .D (n6128),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1290 (
	   .Q (_net_7729),
	   .D (n6124),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1289 (
	   .Q (_net_6181),
	   .D (n6119),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1288 (
	   .Q (net_6804),
	   .D (n6114),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1287 (
	   .Q (net_7372),
	   .D (n6110),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1286 (
	   .Q (net_6686),
	   .D (n6106),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1285 (
	   .Q (net_6763),
	   .D (n6102),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1284 (
	   .Q (net_6335),
	   .D (n6098),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1283 (
	   .Q (_net_7405),
	   .D (n6093),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1282 (
	   .Q (net_6054),
	   .D (n6088),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1281 (
	   .Q (net_261),
	   .D (n6083),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1280 (
	   .Q (_net_7796),
	   .D (n6078),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1279 (
	   .Q (_net_6558),
	   .D (n6074),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1278 (
	   .Q (net_6630),
	   .D (n6069),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1277 (
	   .Q (net_6466),
	   .D (n6066),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1276 (
	   .Q (_net_7482),
	   .D (n6061),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1275 (
	   .Q (net_6802),
	   .D (n6056),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1274 (
	   .Q (_net_6132),
	   .D (n6052),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1273 (
	   .Q (net_6362),
	   .D (n6047),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1272 (
	   .Q (net_6733),
	   .D (n6043),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1271 (
	   .Q (net_251),
	   .D (n6038),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1270 (
	   .Q (net_7125),
	   .D (n6034),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1269 (
	   .Q (_net_6081),
	   .D (n6029),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1268 (
	   .Q (_net_7596),
	   .D (n6024),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1267 (
	   .Q (net_6314),
	   .D (n6019),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1266 (
	   .Q (net_5861),
	   .D (n6014),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1265 (
	   .Q (net_6497),
	   .D (n6009),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1264 (
	   .Q (net_7115),
	   .D (n6006),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1263 (
	   .Q (net_7712),
	   .D (n6002),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1262 (
	   .Q (_net_6066),
	   .D (n5997),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1261 (
	   .Q (_net_7357),
	   .D (n5992),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1260 (
	   .Q (_net_6410),
	   .D (n5987),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1259 (
	   .Q (_net_6689),
	   .D (n5982),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1258 (
	   .Q (net_6618),
	   .D (n5978),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1257 (
	   .Q (_net_7360),
	   .D (n5973),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1256 (
	   .Q (net_7056),
	   .D (n5968),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1255 (
	   .Q (_net_7798),
	   .D (n5964),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1254 (
	   .Q (_net_6006),
	   .D (n5960),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1253 (
	   .Q (net_6255),
	   .D (n5955),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1252 (
	   .Q (net_6973),
	   .D (n5951),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1251 (
	   .Q (net_6562),
	   .D (n5947),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1250 (
	   .Q (net_6887),
	   .D (n5943),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1249 (
	   .Q (_net_7553),
	   .D (n5938),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1248 (
	   .Q (net_7127),
	   .D (n5934),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1247 (
	   .Q (net_6580),
	   .D (n5930),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1246 (
	   .Q (_net_6040),
	   .D (n5925),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1245 (
	   .Q (net_6927),
	   .D (n5920),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1244 (
	   .Q (net_6971),
	   .D (n5917),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1243 (
	   .Q (net_6538),
	   .D (n5912),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1242 (
	   .Q (net_6376),
	   .D (n5908),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1241 (
	   .Q (net_7792),
	   .D (n5903),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1240 (
	   .Q (_net_7407),
	   .D (n5899),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1239 (
	   .Q (net_356),
	   .D (n5894),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1238 (
	   .Q (_net_283),
	   .D (n5890),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1237 (
	   .Q (_net_5982),
	   .D (n5885),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1236 (
	   .Q (net_6720),
	   .D (n5881),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1235 (
	   .Q (net_6954),
	   .D (n5876),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1234 (
	   .Q (net_6340),
	   .D (n5872),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1233 (
	   .Q (net_7306),
	   .D (n5867),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1232 (
	   .Q (net_7102),
	   .D (n5864),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1231 (
	   .Q (net_6479),
	   .D (n5860),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1230 (
	   .Q (net_6416),
	   .D (n5855),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1229 (
	   .Q (_net_7734),
	   .D (n5850),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1228 (
	   .Q (net_259),
	   .D (n5845),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1227 (
	   .Q (net_6925),
	   .D (n5840),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1226 (
	   .Q (net_6934),
	   .D (n5836),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1225 (
	   .Q (net_6878),
	   .D (n5833),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1224 (
	   .Q (net_164),
	   .D (n5828),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1223 (
	   .Q (net_7113),
	   .D (n5824),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1222 (
	   .Q (net_247),
	   .D (n5819),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1221 (
	   .Q (net_7676),
	   .D (n5814),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1220 (
	   .Q (_net_7561),
	   .D (n5809),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1219 (
	   .Q (net_6437),
	   .D (n5805),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1218 (
	   .Q (net_7012),
	   .D (n5801),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1217 (
	   .Q (net_6632),
	   .D (n5796),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1216 (
	   .Q (net_7529),
	   .D (n5792),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1215 (
	   .Q (net_6779),
	   .D (n5787),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1214 (
	   .Q (net_373),
	   .D (n5783),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1213 (
	   .Q (net_6642),
	   .D (n5779),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1212 (
	   .Q (_net_6154),
	   .D (n5775),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1211 (
	   .Q (net_6480),
	   .D (n5771),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1210 (
	   .Q (net_6590),
	   .D (n5767),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1209 (
	   .Q (net_6560),
	   .D (n5763),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1208 (
	   .Q (net_6327),
	   .D (n5758),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1207 (
	   .Q (_net_6414),
	   .D (n5753),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1206 (
	   .Q (_net_6825),
	   .D (n5748),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1205 (
	   .Q (net_7244),
	   .D (n5744),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1204 (
	   .Q (_net_5998),
	   .D (n5739),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1203 (
	   .Q (net_7026),
	   .D (n5735),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1202 (
	   .Q (net_7107),
	   .D (n5731),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1201 (
	   .Q (net_6598),
	   .D (n5727),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1200 (
	   .Q (_net_269),
	   .D (n5722),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1199 (
	   .Q (net_6523),
	   .D (n5717),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1198 (
	   .Q (net_6668),
	   .D (n5713),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1197 (
	   .Q (net_6412),
	   .D (n5709),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1196 (
	   .Q (net_6942),
	   .D (n5704),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1195 (
	   .Q (net_169),
	   .D (n5700),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1194 (
	   .Q (net_6609),
	   .D (n5696),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1193 (
	   .Q (_net_6283),
	   .D (n5691),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l1192 (
	   .Q (_net_7822),
	   .D (n5686),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1191 (
	   .Q (net_7030),
	   .D (n5682),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1190 (
	   .Q (net_6727),
	   .D (n5679),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1189 (
	   .Q (_net_7564),
	   .D (n5674),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1188 (
	   .Q (_net_7380),
	   .D (n5669),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1187 (
	   .Q (net_7215),
	   .D (n5664),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1186 (
	   .Q (net_5849),
	   .D (n5660),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1185 (
	   .Q (net_6490),
	   .D (n5655),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1184 (
	   .Q (net_7202),
	   .D (n5651),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1183 (
	   .Q (net_6983),
	   .D (n5648),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1182 (
	   .Q (_net_7634),
	   .D (n5643),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1181 (
	   .Q (_net_6205),
	   .D (n5638),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1180 (
	   .Q (_net_7736),
	   .D (n5633),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1179 (
	   .Q (net_7647),
	   .D (n5628),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1178 (
	   .Q (_net_6138),
	   .D (n5623),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1177 (
	   .Q (net_6243),
	   .D (n5618),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1176 (
	   .Q (net_7080),
	   .D (n5613),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1175 (
	   .Q (net_133),
	   .D (n5610),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1174 (
	   .Q (net_6368),
	   .D (n5606),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1173 (
	   .Q (_net_7420),
	   .D (n5601),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1172 (
	   .Q (_net_6162),
	   .D (n5596),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1171 (
	   .Q (net_7640),
	   .D (n5591),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1170 (
	   .Q (net_7235),
	   .D (n5588),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1169 (
	   .Q (net_7546),
	   .D (n5584),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1168 (
	   .Q (_net_7622),
	   .D (n5579),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1167 (
	   .Q (net_6620),
	   .D (n5575),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1166 (
	   .Q (_net_7502),
	   .D (n5570),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1165 (
	   .Q (_net_7430),
	   .D (n5565),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1164 (
	   .Q (net_6789),
	   .D (n5560),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1163 (
	   .Q (net_343),
	   .D (n5556),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1162 (
	   .Q (net_7528),
	   .D (n5552),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1161 (
	   .Q (net_6670),
	   .D (n5547),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1160 (
	   .Q (_net_7577),
	   .D (n5543),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1159 (
	   .Q (net_6839),
	   .D (n5539),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1158 (
	   .Q (_net_7721),
	   .D (n5534),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1157 (
	   .Q (net_7780),
	   .D (n5529),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1156 (
	   .Q (x172),
	   .D (n5525),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1155 (
	   .Q (net_7018),
	   .D (n5521),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1154 (
	   .Q (x390),
	   .D (n5517),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1153 (
	   .Q (net_6024),
	   .D (n5513),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1152 (
	   .Q (_net_7467),
	   .D (n5508),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1151 (
	   .Q (net_7100),
	   .D (n5504),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1150 (
	   .Q (net_6575),
	   .D (n5500),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1149 (
	   .Q (_net_270),
	   .D (n5495),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1148 (
	   .Q (_net_7513),
	   .D (n5490),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1147 (
	   .Q (net_390),
	   .D (n5486),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1146 (
	   .Q (net_6915),
	   .D (n5481),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1145 (
	   .Q (_net_7587),
	   .D (n5477),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1144 (
	   .Q (net_7610),
	   .D (n5472),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1143 (
	   .Q (net_6610),
	   .D (n5469),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1142 (
	   .Q (net_7335),
	   .D (n5464),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1141 (
	   .Q (net_6251),
	   .D (n5460),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1140 (
	   .Q (_net_5987),
	   .D (n5455),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1139 (
	   .Q (net_6436),
	   .D (n5451),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1138 (
	   .Q (_net_119),
	   .D (n5446),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1137 (
	   .Q (net_6551),
	   .D (n5441),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1136 (
	   .Q (net_380),
	   .D (n5437),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1135 (
	   .Q (net_6766),
	   .D (n5433),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1134 (
	   .Q (_net_6030),
	   .D (n5429),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1133 (
	   .Q (net_7167),
	   .D (n5424),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1132 (
	   .Q (_net_7295),
	   .D (n5420),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1131 (
	   .Q (net_7206),
	   .D (n5415),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1130 (
	   .Q (_net_7631),
	   .D (n5411),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1129 (
	   .Q (_net_7429),
	   .D (n5406),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1128 (
	   .Q (net_7151),
	   .D (n5402),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1127 (
	   .Q (net_159),
	   .D (n5397),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1126 (
	   .Q (net_7021),
	   .D (n5393),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1125 (
	   .Q (_net_6096),
	   .D (n5388),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1124 (
	   .Q (net_6816),
	   .D (n5383),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1123 (
	   .Q (net_6729),
	   .D (n5380),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1122 (
	   .Q (net_6237),
	   .D (n5375),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1121 (
	   .Q (_net_7657),
	   .D (n5370),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1120 (
	   .Q (net_6860),
	   .D (n5366),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1119 (
	   .Q (net_6460),
	   .D (n5362),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1118 (
	   .Q (net_6454),
	   .D (n5358),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1117 (
	   .Q (_net_7280),
	   .D (n5353),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1116 (
	   .Q (net_6987),
	   .D (n5349),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1115 (
	   .Q (_net_6420),
	   .D (n5344),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1114 (
	   .Q (net_6357),
	   .D (n5339),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1113 (
	   .Q (net_7002),
	   .D (n5335),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1112 (
	   .Q (_net_7662),
	   .D (n5330),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1111 (
	   .Q (net_6844),
	   .D (n5326),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1110 (
	   .Q (_net_7684),
	   .D (n5321),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1109 (
	   .Q (net_6061),
	   .D (n5316),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1108 (
	   .Q (net_7006),
	   .D (n5312),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1107 (
	   .Q (_net_7411),
	   .D (n5307),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1106 (
	   .Q (net_6324),
	   .D (n5302),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1105 (
	   .Q (net_6965),
	   .D (n5298),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1104 (
	   .Q (_net_7599),
	   .D (n5293),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1103 (
	   .Q (net_320),
	   .D (n5288),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1102 (
	   .Q (_net_6284),
	   .D (n5284),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1101 (
	   .Q (_net_7731),
	   .D (n5279),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1100 (
	   .Q (_net_7292),
	   .D (n5274),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1099 (
	   .Q (net_7168),
	   .D (n5269),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1098 (
	   .Q (_net_7416),
	   .D (n5265),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1097 (
	   .Q (net_6843),
	   .D (n5261),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1096 (
	   .Q (_net_7567),
	   .D (n5256),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1095 (
	   .Q (_net_7297),
	   .D (n5251),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1094 (
	   .Q (net_6897),
	   .D (n5246),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1093 (
	   .Q (net_6676),
	   .D (n5242),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1092 (
	   .Q (net_6487),
	   .D (n5239),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1091 (
	   .Q (net_7176),
	   .D (n5234),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1090 (
	   .Q (_net_7422),
	   .D (n5230),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1089 (
	   .Q (_net_7593),
	   .D (n5225),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1088 (
	   .Q (net_6857),
	   .D (n5221),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1087 (
	   .Q (net_6569),
	   .D (n5217),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1086 (
	   .Q (_net_6114),
	   .D (n5212),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1085 (
	   .Q (_net_7686),
	   .D (n5207),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1084 (
	   .Q (net_6506),
	   .D (n5202),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l1083 (
	   .Q (_net_6084),
	   .D (n5198),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1082 (
	   .Q (net_7037),
	   .D (n5193),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1081 (
	   .Q (net_6656),
	   .D (n5189),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1080 (
	   .Q (net_7691),
	   .D (n5186),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1079 (
	   .Q (_net_7803),
	   .D (n5181),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1078 (
	   .Q (net_6841),
	   .D (n5178),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1077 (
	   .Q (net_6940),
	   .D (n5173),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1076 (
	   .Q (_net_7435),
	   .D (n5169),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1075 (
	   .Q (_net_271),
	   .D (n5164),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1074 (
	   .Q (net_130),
	   .D (n5159),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1073 (
	   .Q (net_6428),
	   .D (n5156),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1072 (
	   .Q (net_6516),
	   .D (n5151),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1071 (
	   .Q (net_6572),
	   .D (n5148),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1070 (
	   .Q (_net_7272),
	   .D (n5143),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1069 (
	   .Q (net_6985),
	   .D (n5139),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l1068 (
	   .Q (net_218),
	   .D (n5134),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l1067 (
	   .Q (x149),
	   .D (n5130),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1066 (
	   .Q (net_6589),
	   .D (n5126),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1065 (
	   .Q (net_308),
	   .D (n5121),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1064 (
	   .Q (_net_227),
	   .D (n5117),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1063 (
	   .Q (_net_6415),
	   .D (n5112),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1062 (
	   .Q (net_208),
	   .D (n5107),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1061 (
	   .Q (x379),
	   .D (n5103),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1060 (
	   .Q (net_324),
	   .D (n5098),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1059 (
	   .Q (_net_7433),
	   .D (n5094),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1058 (
	   .Q (net_7011),
	   .D (n5090),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1057 (
	   .Q (net_6057),
	   .D (n5085),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1056 (
	   .Q (_net_7514),
	   .D (n5080),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1055 (
	   .Q (_net_7508),
	   .D (n5075),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1054 (
	   .Q (net_6663),
	   .D (n5070),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1053 (
	   .Q (net_6311),
	   .D (n5066),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1052 (
	   .Q (_net_7507),
	   .D (n5061),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1051 (
	   .Q (net_7376),
	   .D (n5056),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1050 (
	   .Q (net_6970),
	   .D (n5053),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1049 (
	   .Q (net_7614),
	   .D (n5048),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1048 (
	   .Q (net_7399),
	   .D (n5045),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1047 (
	   .Q (_net_6034),
	   .D (n5040),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1046 (
	   .Q (net_7219),
	   .D (n5035),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1045 (
	   .Q (net_6546),
	   .D (n5031),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1044 (
	   .Q (net_7518),
	   .D (n5027),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l1043 (
	   .Q (net_7539),
	   .D (n5023),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1042 (
	   .Q (_net_6693),
	   .D (n5018),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1041 (
	   .Q (_net_7727),
	   .D (n5013),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1040 (
	   .Q (net_331),
	   .D (n5008),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1039 (
	   .Q (net_6854),
	   .D (n5005),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1038 (
	   .Q (net_6617),
	   .D (n5001),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l1037 (
	   .Q (net_6241),
	   .D (n4996),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1036 (
	   .Q (x765),
	   .D (n4992),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l1035 (
	   .Q (_net_7571),
	   .D (n4987),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1034 (
	   .Q (net_6858),
	   .D (n4983),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1033 (
	   .Q (net_6484),
	   .D (n4979),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1032 (
	   .Q (_net_6157),
	   .D (n4974),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1031 (
	   .Q (net_6808),
	   .D (n4969),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l1030 (
	   .Q (net_6923),
	   .D (n4965),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1029 (
	   .Q (_net_7651),
	   .D (n4961),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1028 (
	   .Q (net_6718),
	   .D (n4957),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1027 (
	   .Q (_net_295),
	   .D (n4952),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l1026 (
	   .Q (net_7085),
	   .D (n4947),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1025 (
	   .Q (net_144),
	   .D (n4944),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1024 (
	   .Q (net_7047),
	   .D (n4940),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1023 (
	   .Q (_net_7659),
	   .D (n4936),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l1022 (
	   .Q (net_6820),
	   .D (n4931),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1021 (
	   .Q (_net_7782),
	   .D (n4927),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l1020 (
	   .Q (_net_5970),
	   .D (n4922),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1019 (
	   .Q (_net_6011),
	   .D (n4917),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l1018 (
	   .Q (net_6573),
	   .D (n4913),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l1017 (
	   .Q (_net_5967),
	   .D (n4908),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l1016 (
	   .Q (net_7001),
	   .D (n4904),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1015 (
	   .Q (net_6339),
	   .D (n4899),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l1014 (
	   .Q (net_7154),
	   .D (n4895),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l1013 (
	   .Q (net_7203),
	   .D (n4890),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1012 (
	   .Q (net_202),
	   .D (n4886),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l1011 (
	   .Q (net_349),
	   .D (n4881),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l1010 (
	   .Q (_net_6406),
	   .D (n4877),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l1009 (
	   .Q (_net_284),
	   .D (n4872),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l1008 (
	   .Q (net_7189),
	   .D (n4867),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l1007 (
	   .Q (net_6403),
	   .D (n4862),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1006 (
	   .Q (_net_5975),
	   .D (n4857),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l1005 (
	   .Q (net_6875),
	   .D (n4853),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l1004 (
	   .Q (net_6250),
	   .D (n4848),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1003 (
	   .Q (_net_6019),
	   .D (n4843),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l1002 (
	   .Q (net_6509),
	   .D (n4838),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l1001 (
	   .Q (net_6650),
	   .D (n4834),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l1000 (
	   .Q (x234),
	   .D (n4831),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0999 (
	   .Q (net_6567),
	   .D (n4827),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0998 (
	   .Q (net_7304),
	   .D (n4822),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0997 (
	   .Q (_net_7624),
	   .D (n4818),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0996 (
	   .Q (net_7128),
	   .D (n4814),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0995 (
	   .Q (_net_7655),
	   .D (n4809),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0994 (
	   .Q (net_7014),
	   .D (n4805),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0993 (
	   .Q (_net_7452),
	   .D (n4800),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0992 (
	   .Q (net_6935),
	   .D (n4795),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0991 (
	   .Q (net_6931),
	   .D (n4791),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0990 (
	   .Q (_net_7559),
	   .D (n4787),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0989 (
	   .Q (net_6352),
	   .D (n4782),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0988 (
	   .Q (net_6449),
	   .D (n4778),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0987 (
	   .Q (net_7545),
	   .D (n4774),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0986 (
	   .Q (net_7455),
	   .D (n4769),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0985 (
	   .Q (net_6231),
	   .D (n4765),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0984 (
	   .Q (_net_7706),
	   .D (n4760),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0983 (
	   .Q (net_6349),
	   .D (n4755),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0982 (
	   .Q (net_6334),
	   .D (n4750),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0981 (
	   .Q (net_6502),
	   .D (n4745),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0980 (
	   .Q (net_6735),
	   .D (n4742),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0979 (
	   .Q (_net_7382),
	   .D (n4737),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0978 (
	   .Q (_net_7286),
	   .D (n4732),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0977 (
	   .Q (_net_7692),
	   .D (n4727),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0976 (
	   .Q (net_6271),
	   .D (n4722),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0975 (
	   .Q (net_6544),
	   .D (n4717),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0974 (
	   .Q (net_7142),
	   .D (n4713),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0973 (
	   .Q (_net_6073),
	   .D (n4708),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0972 (
	   .Q (_net_7749),
	   .D (n4703),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0971 (
	   .Q (net_6993),
	   .D (n4699),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0970 (
	   .Q (net_7493),
	   .D (n4694),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0969 (
	   .Q (net_7370),
	   .D (n4690),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0968 (
	   .Q (net_378),
	   .D (n4686),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0967 (
	   .Q (_net_7797),
	   .D (n4681),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0966 (
	   .Q (x744),
	   .D (n4678),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0965 (
	   .Q (net_6055),
	   .D (n4673),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0964 (
	   .Q (net_6581),
	   .D (n4669),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0963 (
	   .Q (net_6736),
	   .D (n4665),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0962 (
	   .Q (net_7197),
	   .D (n4660),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0961 (
	   .Q (_net_7288),
	   .D (n4656),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0960 (
	   .Q (net_6367),
	   .D (n4651),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0959 (
	   .Q (_net_7269),
	   .D (n4646),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0958 (
	   .Q (_net_6064),
	   .D (n4641),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0957 (
	   .Q (net_253),
	   .D (n4636),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0956 (
	   .Q (net_6786),
	   .D (n4631),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0955 (
	   .Q (_net_7346),
	   .D (n4627),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0954 (
	   .Q (net_6273),
	   .D (n4622),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0953 (
	   .Q (net_6637),
	   .D (n4617),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0952 (
	   .Q (net_6776),
	   .D (n4613),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0951 (
	   .Q (_net_7586),
	   .D (n4609),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0950 (
	   .Q (net_6635),
	   .D (n4604),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0949 (
	   .Q (net_7068),
	   .D (n4600),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0948 (
	   .Q (_net_7413),
	   .D (n4596),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0947 (
	   .Q (_net_7233),
	   .D (n4591),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0946 (
	   .Q (_net_6297),
	   .D (n4586),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0945 (
	   .Q (net_7079),
	   .D (n4581),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0944 (
	   .Q (net_6305),
	   .D (n4577),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0943 (
	   .Q (_net_7475),
	   .D (n4572),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0942 (
	   .Q (net_6225),
	   .D (n4567),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0941 (
	   .Q (net_6761),
	   .D (n4562),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0940 (
	   .Q (net_146),
	   .D (n4558),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0939 (
	   .Q (_net_6165),
	   .D (n4553),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0938 (
	   .Q (net_6489),
	   .D (n4548),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0937 (
	   .Q (_net_7480),
	   .D (n4544),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0936 (
	   .Q (_net_6172),
	   .D (n4539),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0935 (
	   .Q (net_6195),
	   .D (n4534),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0934 (
	   .Q (_net_6189),
	   .D (n4529),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0933 (
	   .Q (net_138),
	   .D (n4524),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0932 (
	   .Q (net_246),
	   .D (n4520),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0931 (
	   .Q (_net_6173),
	   .D (n4515),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0930 (
	   .Q (_net_7469),
	   .D (n4510),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0929 (
	   .Q (net_7075),
	   .D (n4505),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0928 (
	   .Q (net_155),
	   .D (n4501),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0927 (
	   .Q (net_389),
	   .D (n4496),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0926 (
	   .Q (_net_6018),
	   .D (n4491),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0925 (
	   .Q (net_7129),
	   .D (n4487),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0924 (
	   .Q (_net_6148),
	   .D (n4482),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0923 (
	   .Q (net_6448),
	   .D (n4478),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0922 (
	   .Q (net_7199),
	   .D (n4473),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0921 (
	   .Q (net_6343),
	   .D (n4469),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0920 (
	   .Q (_net_7323),
	   .D (n4464),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0919 (
	   .Q (net_7741),
	   .D (n4459),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0918 (
	   .Q (x179),
	   .D (n4456),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0917 (
	   .Q (net_7374),
	   .D (n4451),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0916 (
	   .Q (net_6886),
	   .D (n4448),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0915 (
	   .Q (_net_6206),
	   .D (n4443),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0914 (
	   .Q (_net_7403),
	   .D (n4438),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0913 (
	   .Q (_net_7332),
	   .D (n4433),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0912 (
	   .Q (net_7366),
	   .D (n4428),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0911 (
	   .Q (_net_6045),
	   .D (n4424),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0910 (
	   .Q (net_6347),
	   .D (n4419),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0909 (
	   .Q (_net_7718),
	   .D (n4414),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0908 (
	   .Q (net_7111),
	   .D (n4410),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0907 (
	   .Q (_net_265),
	   .D (n4405),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0906 (
	   .Q (net_7162),
	   .D (n4401),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0905 (
	   .Q (net_6564),
	   .D (n4397),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0904 (
	   .Q (_net_7301),
	   .D (n4392),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0903 (
	   .Q (net_6431),
	   .D (n4388),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0902 (
	   .Q (net_6974),
	   .D (n4384),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0901 (
	   .Q (_net_7278),
	   .D (n4379),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0900 (
	   .Q (net_6950),
	   .D (n4374),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0899 (
	   .Q (net_6641),
	   .D (n4370),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0898 (
	   .Q (net_6762),
	   .D (n4365),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0897 (
	   .Q (net_6863),
	   .D (n4362),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0896 (
	   .Q (_net_6009),
	   .D (n4357),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0895 (
	   .Q (net_7646),
	   .D (n4352),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0894 (
	   .Q (_net_7505),
	   .D (n4348),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0893 (
	   .Q (net_7771),
	   .D (n4343),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0892 (
	   .Q (net_6805),
	   .D (n4338),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0891 (
	   .Q (net_7641),
	   .D (n4333),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0890 (
	   .Q (net_6978),
	   .D (n4330),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0889 (
	   .Q (net_6388),
	   .D (n4326),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0888 (
	   .Q (_net_6050),
	   .D (n4322),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0887 (
	   .Q (net_6471),
	   .D (n4318),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0886 (
	   .Q (_net_6422),
	   .D (n4313),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0885 (
	   .Q (net_6753),
	   .D (n4309),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0884 (
	   .Q (_net_7688),
	   .D (n4304),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0883 (
	   .Q (_net_6128),
	   .D (n4299),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0882 (
	   .Q (_net_7318),
	   .D (n4294),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0881 (
	   .Q (_net_229),
	   .D (n4289),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0880 (
	   .Q (_net_7810),
	   .D (n4284),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0879 (
	   .Q (net_6926),
	   .D (n4280),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0878 (
	   .Q (_net_5981),
	   .D (n4276),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0877 (
	   .Q (net_312),
	   .D (n4271),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0876 (
	   .Q (net_7031),
	   .D (n4267),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0875 (
	   .Q (net_7338),
	   .D (n4263),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0874 (
	   .Q (net_296),
	   .D (n4258),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0873 (
	   .Q (net_376),
	   .D (n4253),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0872 (
	   .Q (_net_6152),
	   .D (n4249),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0871 (
	   .Q (net_7398),
	   .D (n4245),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0870 (
	   .Q (_net_7635),
	   .D (n4240),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0869 (
	   .Q (net_6643),
	   .D (n4235),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0868 (
	   .Q (net_5858),
	   .D (n4231),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0867 (
	   .Q (_net_5968),
	   .D (n4226),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0866 (
	   .Q (net_7049),
	   .D (n4221),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0865 (
	   .Q (_net_7630),
	   .D (n4217),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0864 (
	   .Q (net_206),
	   .D (n4212),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0863 (
	   .Q (net_7178),
	   .D (n4207),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0862 (
	   .Q (_net_277),
	   .D (n4203),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0861 (
	   .Q (net_6447),
	   .D (n4199),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0860 (
	   .Q (net_6684),
	   .D (n4194),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0859 (
	   .Q (net_7123),
	   .D (n4191),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0858 (
	   .Q (_net_7321),
	   .D (n4186),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0857 (
	   .Q (net_234),
	   .D (n4181),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0856 (
	   .Q (net_6263),
	   .D (n4176),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0855 (
	   .Q (_net_7784),
	   .D (n4171),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0854 (
	   .Q (_net_7437),
	   .D (n4166),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0853 (
	   .Q (net_367),
	   .D (n4161),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0852 (
	   .Q (net_6714),
	   .D (n4158),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0851 (
	   .Q (_net_6239),
	   .D (n4153),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0850 (
	   .Q (net_7028),
	   .D (n4148),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0849 (
	   .Q (net_6592),
	   .D (n4145),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0848 (
	   .Q (_net_7347),
	   .D (n4140),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0847 (
	   .Q (_net_7232),
	   .D (n4135),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0846 (
	   .Q (net_7400),
	   .D (n4131),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0845 (
	   .Q (_net_7227),
	   .D (n4126),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0844 (
	   .Q (_net_276),
	   .D (n4121),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0843 (
	   .Q (_net_7364),
	   .D (n4116),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0842 (
	   .Q (net_6867),
	   .D (n4112),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0841 (
	   .Q (_net_7719),
	   .D (n4107),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0840 (
	   .Q (net_6778),
	   .D (n4102),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0839 (
	   .Q (net_6493),
	   .D (n4098),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0838 (
	   .Q (_net_7404),
	   .D (n4094),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0837 (
	   .Q (_net_6411),
	   .D (n4089),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0836 (
	   .Q (_net_294),
	   .D (n4084),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0835 (
	   .Q (net_7636),
	   .D (n4079),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0834 (
	   .Q (net_364),
	   .D (n4075),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0833 (
	   .Q (net_6541),
	   .D (n4071),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0832 (
	   .Q (net_6444),
	   .D (n4068),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0831 (
	   .Q (_net_7329),
	   .D (n4063),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0830 (
	   .Q (net_7013),
	   .D (n4059),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0829 (
	   .Q (net_7711),
	   .D (n4055),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0828 (
	   .Q (net_6613),
	   .D (n4051),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0827 (
	   .Q (net_355),
	   .D (n4046),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0826 (
	   .Q (_net_7633),
	   .D (n4042),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0825 (
	   .Q (net_6790),
	   .D (n4037),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0824 (
	   .Q (net_7191),
	   .D (n4033),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0823 (
	   .Q (_net_7601),
	   .D (n4029),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0822 (
	   .Q (net_141),
	   .D (n4024),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0821 (
	   .Q (net_6810),
	   .D (n4020),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0820 (
	   .Q (_net_7733),
	   .D (n4016),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0819 (
	   .Q (net_6279),
	   .D (n4011),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0818 (
	   .Q (net_6852),
	   .D (n4007),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0817 (
	   .Q (net_6949),
	   .D (n4002),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0816 (
	   .Q (_net_7095),
	   .D (n3998),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0815 (
	   .Q (net_7165),
	   .D (n3993),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0814 (
	   .Q (net_309),
	   .D (n3989),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0813 (
	   .Q (net_7050),
	   .D (n3985),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0812 (
	   .Q (_net_6112),
	   .D (n3981),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0811 (
	   .Q (_net_6202),
	   .D (n3976),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0810 (
	   .Q (net_7537),
	   .D (n3972),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0809 (
	   .Q (_net_7510),
	   .D (n3967),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0808 (
	   .Q (net_6372),
	   .D (n3962),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0807 (
	   .Q (net_372),
	   .D (n3957),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0806 (
	   .Q (net_7185),
	   .D (n3953),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0805 (
	   .Q (net_6819),
	   .D (n3949),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0804 (
	   .Q (net_369),
	   .D (n3945),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0803 (
	   .Q (_net_7591),
	   .D (n3941),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0802 (
	   .Q (net_6685),
	   .D (n3936),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0801 (
	   .Q (_net_7418),
	   .D (n3932),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0800 (
	   .Q (_net_7563),
	   .D (n3927),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0799 (
	   .Q (_net_6116),
	   .D (n3922),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0798 (
	   .Q (net_7184),
	   .D (n3917),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0797 (
	   .Q (_net_7270),
	   .D (n3913),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0796 (
	   .Q (net_223),
	   .D (n3908),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0795 (
	   .Q (net_7239),
	   .D (n3904),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0794 (
	   .Q (net_7034),
	   .D (n3899),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0793 (
	   .Q (net_6855),
	   .D (n3896),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0792 (
	   .Q (_net_123),
	   .D (n3891),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0791 (
	   .Q (_net_7574),
	   .D (n3886),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0790 (
	   .Q (net_6899),
	   .D (n3881),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0789 (
	   .Q (_net_6065),
	   .D (n3877),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0788 (
	   .Q (_net_188),
	   .D (n3872),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0787 (
	   .Q (net_6636),
	   .D (n3867),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0786 (
	   .Q (net_6850),
	   .D (n3864),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0785 (
	   .Q (_net_7290),
	   .D (n3859),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0784 (
	   .Q (net_6595),
	   .D (n3855),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0783 (
	   .Q (net_6829),
	   .D (n3851),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0782 (
	   .Q (_net_6158),
	   .D (n3846),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0781 (
	   .Q (_net_7652),
	   .D (n3841),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0780 (
	   .Q (_net_6419),
	   .D (n3836),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0779 (
	   .Q (net_6799),
	   .D (n3831),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0778 (
	   .Q (net_286),
	   .D (n3827),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0777 (
	   .Q (net_6252),
	   .D (n3822),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0776 (
	   .Q (net_339),
	   .D (n3817),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0775 (
	   .Q (net_182),
	   .D (n3813),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0774 (
	   .Q (net_6429),
	   .D (n3809),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0773 (
	   .Q (net_7714),
	   .D (n3805),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0772 (
	   .Q (net_7149),
	   .D (n3801),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0771 (
	   .Q (_net_7785),
	   .D (n3796),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0770 (
	   .Q (net_6666),
	   .D (n3791),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0769 (
	   .Q (_net_7092),
	   .D (n3787),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0768 (
	   .Q (_net_7626),
	   .D (n3782),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0767 (
	   .Q (net_6525),
	   .D (n3777),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0766 (
	   .Q (net_6928),
	   .D (n3773),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0765 (
	   .Q (net_6991),
	   .D (n3770),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0764 (
	   .Q (_net_290),
	   .D (n3765),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0763 (
	   .Q (net_6442),
	   .D (n3761),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0762 (
	   .Q (net_336),
	   .D (n3756),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0761 (
	   .Q (net_6245),
	   .D (n3752),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0760 (
	   .Q (net_6325),
	   .D (n3747),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0759 (
	   .Q (_net_7598),
	   .D (n3742),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0758 (
	   .Q (_net_7444),
	   .D (n3737),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0757 (
	   .Q (net_7799),
	   .D (n3733),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0756 (
	   .Q (net_7048),
	   .D (n3729),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0755 (
	   .Q (net_6881),
	   .D (n3725),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0754 (
	   .Q (net_6268),
	   .D (n3720),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0753 (
	   .Q (net_6486),
	   .D (n3716),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0752 (
	   .Q (net_7775),
	   .D (n3711),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0751 (
	   .Q (net_6721),
	   .D (n3707),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0750 (
	   .Q (net_6976),
	   .D (n3703),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0749 (
	   .Q (_net_5853),
	   .D (n3698),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0748 (
	   .Q (_net_7250),
	   .D (n3693),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0747 (
	   .Q (net_6605),
	   .D (n3689),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0746 (
	   .Q (_net_5854),
	   .D (n3684),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0745 (
	   .Q (net_7171),
	   .D (n3679),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0744 (
	   .Q (_net_7728),
	   .D (n3675),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0743 (
	   .Q (net_7061),
	   .D (n3670),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0742 (
	   .Q (_net_7424),
	   .D (n3666),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0741 (
	   .Q (net_7490),
	   .D (n3661),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0740 (
	   .Q (net_6395),
	   .D (n3658),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0739 (
	   .Q (net_6591),
	   .D (n3655),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0738 (
	   .Q (net_7157),
	   .D (n3651),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0737 (
	   .Q (x217),
	   .D (n3647),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0736 (
	   .Q (net_7737),
	   .D (n3642),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0735 (
	   .Q (net_7378),
	   .D (n3638),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0734 (
	   .Q (_net_7665),
	   .D (n3633),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0733 (
	   .Q (_net_7781),
	   .D (n3628),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0732 (
	   .Q (net_6320),
	   .D (n3623),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0731 (
	   .Q (net_6674),
	   .D (n3618),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0730 (
	   .Q (_net_5988),
	   .D (n3614),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0729 (
	   .Q (_net_6092),
	   .D (n3609),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0728 (
	   .Q (net_7678),
	   .D (n3604),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0727 (
	   .Q (net_6583),
	   .D (n3600),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0726 (
	   .Q (_net_5962),
	   .D (n3595),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0725 (
	   .Q (net_6530),
	   .D (n3590),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0724 (
	   .Q (net_6476),
	   .D (n3587),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0723 (
	   .Q (net_255),
	   .D (n3582),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0722 (
	   .Q (_net_6408),
	   .D (n3577),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0721 (
	   .Q (_net_7703),
	   .D (n3572),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0720 (
	   .Q (net_7672),
	   .D (n3567),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0719 (
	   .Q (net_6873),
	   .D (n3564),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0718 (
	   .Q (net_6505),
	   .D (n3559),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0717 (
	   .Q (net_310),
	   .D (n3555),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0716 (
	   .Q (net_7231),
	   .D (n3551),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0715 (
	   .Q (net_7642),
	   .D (n3546),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0714 (
	   .Q (net_6885),
	   .D (n3542),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0713 (
	   .Q (net_6254),
	   .D (n3537),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0712 (
	   .Q (net_329),
	   .D (n3532),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0711 (
	   .Q (net_7082),
	   .D (n3528),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0710 (
	   .Q (net_6216),
	   .D (n3524),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0709 (
	   .Q (net_6765),
	   .D (n3520),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0708 (
	   .Q (_net_6687),
	   .D (n3516),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0707 (
	   .Q (net_7195),
	   .D (n3511),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0706 (
	   .Q (_net_6078),
	   .D (n3507),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0705 (
	   .Q (net_7766),
	   .D (n3502),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0704 (
	   .Q (net_140),
	   .D (n3497),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0703 (
	   .Q (net_7241),
	   .D (n3494),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0702 (
	   .Q (_net_7362),
	   .D (n3489),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0701 (
	   .Q (_net_6290),
	   .D (n3484),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0700 (
	   .Q (net_6332),
	   .D (n3479),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0699 (
	   .Q (_net_6130),
	   .D (n3474),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0698 (
	   .Q (net_7213),
	   .D (n3469),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0697 (
	   .Q (_net_191),
	   .D (n3464),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0696 (
	   .Q (_net_6075),
	   .D (n3459),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0695 (
	   .Q (x786),
	   .D (n3455),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0694 (
	   .Q (net_6369),
	   .D (n3450),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0693 (
	   .Q (net_334),
	   .D (n3445),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0692 (
	   .Q (_net_211),
	   .D (n3440),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0691 (
	   .Q (net_7120),
	   .D (n3436),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0690 (
	   .Q (net_7743),
	   .D (n3431),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0689 (
	   .Q (_net_7618),
	   .D (n3427),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0688 (
	   .Q (net_197),
	   .D (n3422),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0687 (
	   .Q (net_7248),
	   .D (n3418),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0686 (
	   .Q (net_6214),
	   .D (n3413),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0685 (
	   .Q (net_6547),
	   .D (n3408),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0684 (
	   .Q (net_371),
	   .D (n3404),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0683 (
	   .Q (_net_7619),
	   .D (n3400),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0682 (
	   .Q (_net_6142),
	   .D (n3395),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0681 (
	   .Q (_net_7814),
	   .D (n3390),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0680 (
	   .Q (net_7042),
	   .D (n3386),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0679 (
	   .Q (net_6485),
	   .D (n3383),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0678 (
	   .Q (net_6698),
	   .D (n3379),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0677 (
	   .Q (net_7517),
	   .D (n3374),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0676 (
	   .Q (_net_5980),
	   .D (n3370),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0675 (
	   .Q (net_6548),
	   .D (n3365),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0674 (
	   .Q (net_6247),
	   .D (n3361),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0673 (
	   .Q (_net_7583),
	   .D (n3356),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0672 (
	   .Q (x589),
	   .D (n3352),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0671 (
	   .Q (net_7140),
	   .D (n3348),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0670 (
	   .Q (_net_6199),
	   .D (n3343),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0669 (
	   .Q (_net_6041),
	   .D (n3338),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0668 (
	   .Q (net_7344),
	   .D (n3333),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0667 (
	   .Q (net_6868),
	   .D (n3330),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0666 (
	   .Q (net_7310),
	   .D (n3325),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0665 (
	   .Q (x447),
	   .D (n3322),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0664 (
	   .Q (net_6883),
	   .D (n3318),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0663 (
	   .Q (_net_6171),
	   .D (n3313),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0662 (
	   .Q (_net_7266),
	   .D (n3308),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0661 (
	   .Q (net_6536),
	   .D (n3303),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0660 (
	   .Q (net_6623),
	   .D (n3299),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0659 (
	   .Q (_net_6083),
	   .D (n3294),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0658 (
	   .Q (net_7710),
	   .D (n3290),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0657 (
	   .Q (_net_6204),
	   .D (n3285),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0656 (
	   .Q (net_6760),
	   .D (n3280),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0655 (
	   .Q (net_7488),
	   .D (n3276),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0654 (
	   .Q (net_6661),
	   .D (n3272),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0653 (
	   .Q (_net_6102),
	   .D (n3268),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0652 (
	   .Q (_net_116),
	   .D (n3263),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0651 (
	   .Q (_net_7821),
	   .D (n3258),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0650 (
	   .Q (_net_272),
	   .D (n3254),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0649 (
	   .Q (_net_6259),
	   .D (n3249),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0648 (
	   .Q (net_6652),
	   .D (n3244),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0647 (
	   .Q (_net_6175),
	   .D (n3240),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0646 (
	   .Q (_net_7812),
	   .D (n3235),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0645 (
	   .Q (_net_154),
	   .D (n3231),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0644 (
	   .Q (net_6233),
	   .D (n3226),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0643 (
	   .Q (_net_7478),
	   .D (n3222),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0642 (
	   .Q (_net_6110),
	   .D (n3217),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0641 (
	   .Q (_net_7326),
	   .D (n3212),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0640 (
	   .Q (net_6488),
	   .D (n3207),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0639 (
	   .Q (_net_178),
	   .D (n3203),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0638 (
	   .Q (net_7536),
	   .D (n3199),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0637 (
	   .Q (_net_7277),
	   .D (n3194),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0636 (
	   .Q (net_6861),
	   .D (n3190),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0635 (
	   .Q (net_135),
	   .D (n3186),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0634 (
	   .Q (_net_7350),
	   .D (n3182),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0633 (
	   .Q (net_6450),
	   .D (n3178),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0632 (
	   .Q (net_152),
	   .D (n3174),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0631 (
	   .Q (_net_7470),
	   .D (n3170),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0630 (
	   .Q (net_7738),
	   .D (n3165),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0629 (
	   .Q (net_6751),
	   .D (n3162),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0628 (
	   .Q (_net_7690),
	   .D (n3157),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0627 (
	   .Q (net_7040),
	   .D (n3152),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0626 (
	   .Q (_net_7449),
	   .D (n3148),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0625 (
	   .Q (net_6681),
	   .D (n3143),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0624 (
	   .Q (_net_7557),
	   .D (n3139),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0623 (
	   .Q (net_6639),
	   .D (n3134),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0622 (
	   .Q (_net_7410),
	   .D (n3130),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0621 (
	   .Q (net_7387),
	   .D (n3126),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0620 (
	   .Q (net_7643),
	   .D (n3121),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0619 (
	   .Q (net_153),
	   .D (n3117),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0618 (
	   .Q (net_6743),
	   .D (n3114),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0617 (
	   .Q (net_6473),
	   .D (n3110),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0616 (
	   .Q (net_303),
	   .D (n3105),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0615 (
	   .Q (net_6706),
	   .D (n3102),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0614 (
	   .Q (_net_128),
	   .D (n3097),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0613 (
	   .Q (_net_6281),
	   .D (n3092),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0612 (
	   .Q (_net_6688),
	   .D (n3087),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0611 (
	   .Q (net_6796),
	   .D (n3082),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0610 (
	   .Q (net_233),
	   .D (n3078),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0609 (
	   .Q (net_6717),
	   .D (n3074),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0608 (
	   .Q (net_6938),
	   .D (n3069),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0607 (
	   .Q (_net_184),
	   .D (n3065),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0606 (
	   .Q (net_7121),
	   .D (n3061),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0605 (
	   .Q (_net_226),
	   .D (n3056),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0604 (
	   .Q (net_7136),
	   .D (n3052),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0603 (
	   .Q (_net_7667),
	   .D (n3047),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0602 (
	   .Q (_net_6023),
	   .D (n3042),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0601 (
	   .Q (net_6909),
	   .D (n3037),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0600 (
	   .Q (net_6906),
	   .D (n3033),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0599 (
	   .Q (net_7105),
	   .D (n3030),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0598 (
	   .Q (_net_173),
	   .D (n3025),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0597 (
	   .Q (_net_7320),
	   .D (n3020),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0596 (
	   .Q (net_7609),
	   .D (n3015),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0595 (
	   .Q (_net_7751),
	   .D (n3010),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0594 (
	   .Q (_net_6090),
	   .D (n3005),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0593 (
	   .Q (_net_6038),
	   .D (n3000),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0592 (
	   .Q (net_6438),
	   .D (n2996),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0591 (
	   .Q (_net_7531),
	   .D (n2991),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0590 (
	   .Q (_net_6063),
	   .D (n2986),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0589 (
	   .Q (_net_6553),
	   .D (n2981),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0588 (
	   .Q (_net_266),
	   .D (n2976),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0587 (
	   .Q (net_7007),
	   .D (n2972),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0586 (
	   .Q (net_337),
	   .D (n2967),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0585 (
	   .Q (net_6338),
	   .D (n2963),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0584 (
	   .Q (net_7457),
	   .D (n2958),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0583 (
	   .Q (_net_7552),
	   .D (n2953),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0582 (
	   .Q (_net_5969),
	   .D (n2948),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0581 (
	   .Q (net_7158),
	   .D (n2944),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0580 (
	   .Q (net_6781),
	   .D (n2939),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0579 (
	   .Q (_net_5920),
	   .D (n2935),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0578 (
	   .Q (_net_6221),
	   .D (n2930),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0577 (
	   .Q (net_6755),
	   .D (n2926),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0576 (
	   .Q (net_7022),
	   .D (n2922),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0575 (
	   .Q (x315),
	   .D (n2918),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0574 (
	   .Q (net_7336),
	   .D (n2913),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0573 (
	   .Q (net_6946),
	   .D (n2908),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0572 (
	   .Q (net_7461),
	   .D (n2904),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0571 (
	   .Q (_net_7722),
	   .D (n2900),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0570 (
	   .Q (net_7756),
	   .D (n2895),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0569 (
	   .Q (_net_7572),
	   .D (n2890),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0568 (
	   .Q (net_6813),
	   .D (n2885),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0567 (
	   .Q (net_7547),
	   .D (n2882),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0566 (
	   .Q (net_6244),
	   .D (n2877),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0565 (
	   .Q (net_6578),
	   .D (n2873),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0564 (
	   .Q (net_6478),
	   .D (n2869),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0563 (
	   .Q (net_6246),
	   .D (n2864),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0562 (
	   .Q (net_7236),
	   .D (n2860),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0561 (
	   .Q (_net_7501),
	   .D (n2855),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0560 (
	   .Q (net_7670),
	   .D (n2850),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0559 (
	   .Q (_net_7261),
	   .D (n2845),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0558 (
	   .Q (net_6631),
	   .D (n2840),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0557 (
	   .Q (_net_6029),
	   .D (n2836),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0556 (
	   .Q (_net_6156),
	   .D (n2831),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0555 (
	   .Q (net_7153),
	   .D (n2827),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0554 (
	   .Q (net_7024),
	   .D (n2823),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0553 (
	   .Q (net_6579),
	   .D (n2819),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0552 (
	   .Q (net_6539),
	   .D (n2814),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0551 (
	   .Q (_net_214),
	   .D (n2810),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0550 (
	   .Q (_net_7820),
	   .D (n2805),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0549 (
	   .Q (net_6524),
	   .D (n2801),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0548 (
	   .Q (net_232),
	   .D (n2797),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0547 (
	   .Q (net_6664),
	   .D (n2792),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0546 (
	   .Q (net_6496),
	   .D (n2788),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0545 (
	   .Q (net_7343),
	   .D (n2784),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0544 (
	   .Q (net_6880),
	   .D (n2781),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0543 (
	   .Q (_net_5978),
	   .D (n2776),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0542 (
	   .Q (_net_6022),
	   .D (n2771),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0541 (
	   .Q (net_7108),
	   .D (n2767),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0540 (
	   .Q (net_7225),
	   .D (n2762),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0539 (
	   .Q (_net_6097),
	   .D (n2758),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0538 (
	   .Q (net_163),
	   .D (n2753),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0537 (
	   .Q (net_6955),
	   .D (n2748),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0536 (
	   .Q (net_6725),
	   .D (n2745),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0535 (
	   .Q (net_6586),
	   .D (n2741),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0534 (
	   .Q (net_7708),
	   .D (n2737),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0533 (
	   .Q (_net_7314),
	   .D (n2732),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0532 (
	   .Q (net_346),
	   .D (n2727),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0531 (
	   .Q (_net_280),
	   .D (n2723),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0530 (
	   .Q (net_238),
	   .D (n2718),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0529 (
	   .Q (_net_126),
	   .D (n2713),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0528 (
	   .Q (net_6969),
	   .D (n2709),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0527 (
	   .Q (net_6434),
	   .D (n2705),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0526 (
	   .Q (net_6981),
	   .D (n2701),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0525 (
	   .Q (_net_6822),
	   .D (n2696),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0524 (
	   .Q (net_7393),
	   .D (n2692),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0523 (
	   .Q (net_7777),
	   .D (n2687),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0522 (
	   .Q (net_7057),
	   .D (n2682),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0521 (
	   .Q (net_6964),
	   .D (n2679),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0520 (
	   .Q (net_6890),
	   .D (n2675),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0519 (
	   .Q (net_6330),
	   .D (n2670),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0518 (
	   .Q (_net_6121),
	   .D (n2665),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0517 (
	   .Q (net_6215),
	   .D (n2660),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0516 (
	   .Q (net_6606),
	   .D (n2656),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0515 (
	   .Q (net_187),
	   .D (n2651),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0514 (
	   .Q (net_6588),
	   .D (n2647),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0513 (
	   .Q (net_6341),
	   .D (n2642),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0512 (
	   .Q (net_257),
	   .D (n2637),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0511 (
	   .Q (_net_7765),
	   .D (n2632),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0510 (
	   .Q (net_6322),
	   .D (n2627),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0509 (
	   .Q (net_7089),
	   .D (n2622),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0508 (
	   .Q (net_7060),
	   .D (n2618),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0507 (
	   .Q (net_6967),
	   .D (n2615),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0506 (
	   .Q (net_6377),
	   .D (n2610),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0505 (
	   .Q (net_6513),
	   .D (n2605),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0504 (
	   .Q (net_6517),
	   .D (n2601),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0503 (
	   .Q (net_7032),
	   .D (n2597),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0502 (
	   .Q (net_6391),
	   .D (n2594),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0501 (
	   .Q (net_7096),
	   .D (n2590),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0500 (
	   .Q (net_7779),
	   .D (n2585),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0499 (
	   .Q (net_207),
	   .D (n2580),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0498 (
	   .Q (_net_176),
	   .D (n2575),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0497 (
	   .Q (net_6898),
	   .D (n2570),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0496 (
	   .Q (_net_7663),
	   .D (n2566),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0495 (
	   .Q (net_300),
	   .D (n2561),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0494 (
	   .Q (net_6951),
	   .D (n2556),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0493 (
	   .Q (_net_7445),
	   .D (n2552),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0492 (
	   .Q (net_7337),
	   .D (n2547),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0491 (
	   .Q (net_6939),
	   .D (n2543),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0490 (
	   .Q (net_134),
	   .D (n2539),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0489 (
	   .Q (_net_6160),
	   .D (n2534),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0488 (
	   .Q (_net_7419),
	   .D (n2529),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0487 (
	   .Q (net_179),
	   .D (n2524),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0486 (
	   .Q (net_6522),
	   .D (n2519),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0485 (
	   .Q (net_6014),
	   .D (n2515),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0484 (
	   .Q (net_252),
	   .D (n2510),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0483 (
	   .Q (_net_7704),
	   .D (n2505),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0482 (
	   .Q (net_7639),
	   .D (n2500),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0481 (
	   .Q (net_7207),
	   .D (n2496),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0480 (
	   .Q (net_6435),
	   .D (n2493),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0479 (
	   .Q (net_6764),
	   .D (n2488),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0478 (
	   .Q (net_224),
	   .D (n2484),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0477 (
	   .Q (_net_7294),
	   .D (n2479),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0476 (
	   .Q (net_6672),
	   .D (n2474),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0475 (
	   .Q (_net_6118),
	   .D (n2470),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0474 (
	   .Q (net_6918),
	   .D (n2465),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0473 (
	   .Q (net_6426),
	   .D (n2462),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0472 (
	   .Q (_net_5984),
	   .D (n2457),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0471 (
	   .Q (net_6821),
	   .D (n2452),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0470 (
	   .Q (net_377),
	   .D (n2448),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0469 (
	   .Q (_net_5972),
	   .D (n2444),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0468 (
	   .Q (net_7240),
	   .D (n2440),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0467 (
	   .Q (_net_279),
	   .D (n2435),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0466 (
	   .Q (_net_7431),
	   .D (n2430),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0465 (
	   .Q (net_6833),
	   .D (n2426),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0464 (
	   .Q (net_7016),
	   .D (n2422),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0463 (
	   .Q (net_6680),
	   .D (n2417),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0462 (
	   .Q (x699),
	   .D (n2414),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0461 (
	   .Q (_net_7511),
	   .D (n2409),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0460 (
	   .Q (net_7608),
	   .D (n2404),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0459 (
	   .Q (net_6758),
	   .D (n2399),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0458 (
	   .Q (net_183),
	   .D (n2395),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0457 (
	   .Q (net_6576),
	   .D (n2391),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0456 (
	   .Q (_net_6169),
	   .D (n2386),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0455 (
	   .Q (net_7527),
	   .D (n2381),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0454 (
	   .Q (_net_7720),
	   .D (n2377),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0453 (
	   .Q (net_6398),
	   .D (n2373),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0452 (
	   .Q (net_6593),
	   .D (n2370),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0451 (
	   .Q (_net_6163),
	   .D (n2365),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0450 (
	   .Q (net_6912),
	   .D (n2360),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0449 (
	   .Q (net_6277),
	   .D (n2355),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0448 (
	   .Q (net_6236),
	   .D (n2350),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0447 (
	   .Q (net_6849),
	   .D (n2347),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0446 (
	   .Q (net_6501),
	   .D (n2342),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0445 (
	   .Q (net_6920),
	   .D (n2338),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0444 (
	   .Q (_net_7747),
	   .D (n2334),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0443 (
	   .Q (_net_6134),
	   .D (n2329),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0442 (
	   .Q (net_323),
	   .D (n2324),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0441 (
	   .Q (net_7159),
	   .D (n2321),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0440 (
	   .Q (net_6035),
	   .D (n2316),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0439 (
	   .Q (_net_7556),
	   .D (n2312),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0438 (
	   .Q (net_7194),
	   .D (n2307),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0437 (
	   .Q (_net_6187),
	   .D (n2303),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0436 (
	   .Q (_net_6015),
	   .D (n2298),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0435 (
	   .Q (net_6366),
	   .D (n2293),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0434 (
	   .Q (net_142),
	   .D (n2288),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0433 (
	   .Q (net_322),
	   .D (n2284),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0432 (
	   .Q (_net_7748),
	   .D (n2280),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0431 (
	   .Q (_net_6139),
	   .D (n2275),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0430 (
	   .Q (_net_5977),
	   .D (n2270),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0429 (
	   .Q (_net_7401),
	   .D (n2265),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0428 (
	   .Q (net_7671),
	   .D (n2260),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0427 (
	   .Q (net_7458),
	   .D (n2256),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0426 (
	   .Q (_net_6401),
	   .D (n2251),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0425 (
	   .Q (x494),
	   .D (n2247),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0424 (
	   .Q (_net_7724),
	   .D (n2242),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0423 (
	   .Q (_net_6184),
	   .D (n2237),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0422 (
	   .Q (_net_263),
	   .D (n2232),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0421 (
	   .Q (_net_6960),
	   .D (n2227),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0420 (
	   .Q (net_6556),
	   .D (n2222),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0419 (
	   .Q (net_6456),
	   .D (n2218),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0418 (
	   .Q (_net_6016),
	   .D (n2213),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0417 (
	   .Q (_net_5963),
	   .D (n2208),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0416 (
	   .Q (net_6658),
	   .D (n2203),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0415 (
	   .Q (_net_7229),
	   .D (n2199),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0414 (
	   .Q (_net_6177),
	   .D (n2194),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0413 (
	   .Q (net_6540),
	   .D (n2189),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0412 (
	   .Q (net_6443),
	   .D (n2186),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0411 (
	   .Q (_net_7763),
	   .D (n2181),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0410 (
	   .Q (x397),
	   .D (n2177),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0409 (
	   .Q (_net_6963),
	   .D (n2172),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0408 (
	   .Q (_net_7649),
	   .D (n2167),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0407 (
	   .Q (_net_7554),
	   .D (n2162),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0406 (
	   .Q (net_6336),
	   .D (n2157),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0405 (
	   .Q (net_7613),
	   .D (n2152),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0404 (
	   .Q (net_7144),
	   .D (n2149),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0403 (
	   .Q (net_7179),
	   .D (n2144),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0402 (
	   .Q (_net_7683),
	   .D (n2140),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0401 (
	   .Q (net_6730),
	   .D (n2136),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0400 (
	   .Q (net_7147),
	   .D (n2132),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0399 (
	   .Q (net_6310),
	   .D (n2127),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0398 (
	   .Q (net_7076),
	   .D (n2122),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0397 (
	   .Q (net_6603),
	   .D (n2119),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0396 (
	   .Q (net_6452),
	   .D (n2115),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0395 (
	   .Q (net_7003),
	   .D (n2111),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0394 (
	   .Q (net_6191),
	   .D (n2106),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0393 (
	   .Q (net_6741),
	   .D (n2102),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0392 (
	   .Q (net_6709),
	   .D (n2098),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0391 (
	   .Q (net_6893),
	   .D (n2093),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0390 (
	   .Q (net_7063),
	   .D (n2088),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0389 (
	   .Q (net_7371),
	   .D (n2084),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0388 (
	   .Q (net_7754),
	   .D (n2079),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0387 (
	   .Q (net_7201),
	   .D (n2074),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0386 (
	   .Q (_net_6827),
	   .D (n2070),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0385 (
	   .Q (_net_6125),
	   .D (n2065),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0384 (
	   .Q (_net_7352),
	   .D (n2060),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0383 (
	   .Q (_net_7465),
	   .D (n2055),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0382 (
	   .Q (net_7391),
	   .D (n2051),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0381 (
	   .Q (_net_7093),
	   .D (n2046),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0380 (
	   .Q (_net_7483),
	   .D (n2041),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0379 (
	   .Q (net_319),
	   .D (n2036),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0378 (
	   .Q (net_6318),
	   .D (n2031),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0377 (
	   .Q (_net_6107),
	   .D (n2026),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0376 (
	   .Q (net_7790),
	   .D (n2021),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0375 (
	   .Q (_net_7426),
	   .D (n2016),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0374 (
	   .Q (net_7188),
	   .D (n2011),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0373 (
	   .Q (net_6812),
	   .D (n2007),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0372 (
	   .Q (net_6303),
	   .D (n2002),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0371 (
	   .Q (net_6737),
	   .D (n1998),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0370 (
	   .Q (net_7520),
	   .D (n1993),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0369 (
	   .Q (_net_6108),
	   .D (n1988),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0368 (
	   .Q (net_6274),
	   .D (n1983),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0367 (
	   .Q (net_7174),
	   .D (n1978),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0366 (
	   .Q (net_6800),
	   .D (n1973),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0365 (
	   .Q (_net_7594),
	   .D (n1969),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0364 (
	   .Q (net_6346),
	   .D (n1964),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0363 (
	   .Q (_net_129),
	   .D (n1959),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0362 (
	   .Q (net_7052),
	   .D (n1954),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0361 (
	   .Q (_net_7532),
	   .D (n1950),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0360 (
	   .Q (_net_7472),
	   .D (n1945),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0359 (
	   .Q (net_6433),
	   .D (n1941),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0358 (
	   .Q (net_241),
	   .D (n1936),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0357 (
	   .Q (net_6995),
	   .D (n1932),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0356 (
	   .Q (_net_6690),
	   .D (n1927),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0355 (
	   .Q (_net_6070),
	   .D (n1922),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0354 (
	   .Q (net_7116),
	   .D (n1918),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0353 (
	   .Q (net_6543),
	   .D (n1913),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0352 (
	   .Q (_net_7379),
	   .D (n1908),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0351 (
	   .Q (net_6258),
	   .D (n1903),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0350 (
	   .Q (net_6053),
	   .D (n1898),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0349 (
	   .Q (_net_6155),
	   .D (n1893),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0348 (
	   .Q (_net_7628),
	   .D (n1888),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0347 (
	   .Q (_net_6067),
	   .D (n1883),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0346 (
	   .Q (_net_7600),
	   .D (n1878),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0345 (
	   .Q (net_6599),
	   .D (n1874),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0344 (
	   .Q (_net_7255),
	   .D (n1869),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0343 (
	   .Q (net_6699),
	   .D (n1865),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0342 (
	   .Q (net_7767),
	   .D (n1860),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0341 (
	   .Q (_net_7819),
	   .D (n1855),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0340 (
	   .Q (net_6223),
	   .D (n1851),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0339 (
	   .Q (_net_6292),
	   .D (n1846),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0338 (
	   .Q (_net_6087),
	   .D (n1841),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0337 (
	   .Q (_net_7813),
	   .D (n1836),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0336 (
	   .Q (_net_7650),
	   .D (n1832),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0335 (
	   .Q (net_6248),
	   .D (n1827),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0334 (
	   .Q (net_6269),
	   .D (n1822),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0333 (
	   .Q (net_6371),
	   .D (n1817),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0332 (
	   .Q (_net_7359),
	   .D (n1812),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0331 (
	   .Q (_net_7328),
	   .D (n1807),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0330 (
	   .Q (_net_6185),
	   .D (n1802),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0329 (
	   .Q (net_6316),
	   .D (n1797),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0328 (
	   .Q (net_7742),
	   .D (n1792),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0327 (
	   .Q (_net_6296),
	   .D (n1787),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0326 (
	   .Q (net_7035),
	   .D (n1782),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0325 (
	   .Q (net_7551),
	   .D (n1779),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0324 (
	   .Q (net_6602),
	   .D (n1775),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0323 (
	   .Q (_net_5985),
	   .D (n1770),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0322 (
	   .Q (net_7223),
	   .D (n1765),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0321 (
	   .Q (net_6570),
	   .D (n1761),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0320 (
	   .Q (net_6896),
	   .D (n1756),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0319 (
	   .Q (net_7495),
	   .D (n1752),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0318 (
	   .Q (_net_6077),
	   .D (n1747),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0317 (
	   .Q (_net_5996),
	   .D (n1742),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0316 (
	   .Q (_net_7468),
	   .D (n1737),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0315 (
	   .Q (net_6806),
	   .D (n1732),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0314 (
	   .Q (_net_6180),
	   .D (n1727),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0313 (
	   .Q (net_7220),
	   .D (n1722),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0312 (
	   .Q (net_6903),
	   .D (n1718),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0311 (
	   .Q (_net_7358),
	   .D (n1714),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0310 (
	   .Q (net_7170),
	   .D (n1709),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0309 (
	   .Q (net_6500),
	   .D (n1704),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0308 (
	   .Q (net_6432),
	   .D (n1701),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0307 (
	   .Q (_net_6168),
	   .D (n1696),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0306 (
	   .Q (net_6770),
	   .D (n1691),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0305 (
	   .Q (net_6512),
	   .D (n1686),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0304 (
	   .Q (net_6654),
	   .D (n1681),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0303 (
	   .Q (_net_6042),
	   .D (n1677),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0302 (
	   .Q (net_6723),
	   .D (n1673),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0301 (
	   .Q (net_7760),
	   .D (n1668),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0300 (
	   .Q (net_6197),
	   .D (n1663),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0299 (
	   .Q (net_245),
	   .D (n1658),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0298 (
	   .Q (net_6229),
	   .D (n1653),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0297 (
	   .Q (net_7124),
	   .D (n1649),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0296 (
	   .Q (net_260),
	   .D (n1644),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0295 (
	   .Q (net_7308),
	   .D (n1639),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0294 (
	   .Q (_net_7570),
	   .D (n1634),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0293 (
	   .Q (net_6537),
	   .D (n1629),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0292 (
	   .Q (_net_7696),
	   .D (n1624),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0291 (
	   .Q (net_7198),
	   .D (n1619),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0290 (
	   .Q (net_6914),
	   .D (n1615),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0289 (
	   .Q (_net_7498),
	   .D (n1610),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0288 (
	   .Q (net_165),
	   .D (n1605),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0287 (
	   .Q (_net_7759),
	   .D (n1600),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0286 (
	   .Q (net_6732),
	   .D (n1596),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0285 (
	   .Q (net_352),
	   .D (n1591),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0284 (
	   .Q (net_6584),
	   .D (n1587),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0283 (
	   .Q (_net_7535),
	   .D (n1582),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0282 (
	   .Q (net_353),
	   .D (n1577),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0281 (
	   .Q (net_258),
	   .D (n1572),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0280 (
	   .Q (net_6888),
	   .D (n1568),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0279 (
	   .Q (net_6482),
	   .D (n1564),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0278 (
	   .Q (net_7126),
	   .D (n1560),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0277 (
	   .Q (_net_7406),
	   .D (n1555),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0276 (
	   .Q (net_7146),
	   .D (n1551),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0275 (
	   .Q (_net_7534),
	   .D (n1546),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0274 (
	   .Q (x287),
	   .D (n1542),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0273 (
	   .Q (net_7247),
	   .D (n1538),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0272 (
	   .Q (net_203),
	   .D (n1533),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0271 (
	   .Q (net_6375),
	   .D (n1528),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0270 (
	   .Q (net_7106),
	   .D (n1524),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0269 (
	   .Q (_net_6095),
	   .D (n1519),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0268 (
	   .Q (net_6619),
	   .D (n1515),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0267 (
	   .Q (net_7091),
	   .D (n1510),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0266 (
	   .Q (net_7550),
	   .D (n1506),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0265 (
	   .Q (_net_7698),
	   .D (n1501),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0264 (
	   .Q (net_6059),
	   .D (n1496),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0263 (
	   .Q (net_6768),
	   .D (n1491),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0262 (
	   .Q (_net_7746),
	   .D (n1487),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0261 (
	   .Q (_net_7815),
	   .D (n1482),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0260 (
	   .Q (net_6302),
	   .D (n1478),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0259 (
	   .Q (net_6612),
	   .D (n1474),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0258 (
	   .Q (net_357),
	   .D (n1469),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0257 (
	   .Q (net_6953),
	   .D (n1465),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0256 (
	   .Q (net_6328),
	   .D (n1460),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0255 (
	   .Q (net_6633),
	   .D (n1455),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0254 (
	   .Q (_net_6044),
	   .D (n1451),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0253 (
	   .Q (net_6913),
	   .D (n1446),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0252 (
	   .Q (_net_7565),
	   .D (n1442),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0251 (
	   .Q (net_6745),
	   .D (n1438),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0250 (
	   .Q (_net_7768),
	   .D (n1433),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0249 (
	   .Q (_net_7497),
	   .D (n1428),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0248 (
	   .Q (net_6941),
	   .D (n1423),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0247 (
	   .Q (_net_7253),
	   .D (n1419),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0246 (
	   .Q (net_7217),
	   .D (n1414),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0245 (
	   .Q (_net_5960),
	   .D (n1410),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0244 (
	   .Q (_net_6182),
	   .D (n1405),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0243 (
	   .Q (net_6624),
	   .D (n1400),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0242 (
	   .Q (net_6190),
	   .D (n1396),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0241 (
	   .Q (_net_7658),
	   .D (n1391),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0240 (
	   .Q (net_325),
	   .D (n1386),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0239 (
	   .Q (net_6694),
	   .D (n1383),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0238 (
	   .Q (net_7750),
	   .D (n1378),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0237 (
	   .Q (_net_5997),
	   .D (n1373),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0236 (
	   .Q (net_6025),
	   .D (n1368),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0235 (
	   .Q (_net_213),
	   .D (n1363),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0234 (
	   .Q (net_7234),
	   .D (n1359),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0233 (
	   .Q (net_6877),
	   .D (n1355),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0232 (
	   .Q (net_7303),
	   .D (n1350),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0231 (
	   .Q (net_6961),
	   .D (n1345),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0230 (
	   .Q (_net_7707),
	   .D (n1340),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0229 (
	   .Q (_net_5991),
	   .D (n1335),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0228 (
	   .Q (net_6859),
	   .D (n1331),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0227 (
	   .Q (net_6515),
	   .D (n1326),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0226 (
	   .Q (net_7200),
	   .D (n1322),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0225 (
	   .Q (net_7182),
	   .D (n1318),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0224 (
	   .Q (_net_6000),
	   .D (n1314),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0223 (
	   .Q (_net_5966),
	   .D (n1309),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0222 (
	   .Q (net_7395),
	   .D (n1305),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0221 (
	   .Q (net_7070),
	   .D (n1300),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0220 (
	   .Q (_net_7315),
	   .D (n1295),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0219 (
	   .Q (net_6574),
	   .D (n1291),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0218 (
	   .Q (net_7119),
	   .D (n1287),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0217 (
	   .Q (_net_299),
	   .D (n1282),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0216 (
	   .Q (net_7453),
	   .D (n1277),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0215 (
	   .Q (_net_273),
	   .D (n1272),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0214 (
	   .Q (_net_7590),
	   .D (n1267),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0213 (
	   .Q (net_6354),
	   .D (n1262),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0212 (
	   .Q (net_7019),
	   .D (n1258),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0211 (
	   .Q (_net_7512),
	   .D (n1253),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0210 (
	   .Q (net_6759),
	   .D (n1248),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0209 (
	   .Q (net_360),
	   .D (n1244),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0208 (
	   .Q (net_6952),
	   .D (n1240),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0207 (
	   .Q (net_7675),
	   .D (n1236),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0206 (
	   .Q (net_132),
	   .D (n1232),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0205 (
	   .Q (_net_7730),
	   .D (n1228),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0204 (
	   .Q (net_6608),
	   .D (n1224),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0203 (
	   .Q (_net_7428),
	   .D (n1219),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0202 (
	   .Q (_net_7503),
	   .D (n1214),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0201 (
	   .Q (net_6845),
	   .D (n1210),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0200 (
	   .Q (net_7081),
	   .D (n1205),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0199 (
	   .Q (net_6240),
	   .D (n1200),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0198 (
	   .Q (net_6922),
	   .D (n1195),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0197 (
	   .Q (net_6788),
	   .D (n1191),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0196 (
	   .Q (net_345),
	   .D (n1187),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0195 (
	   .Q (net_6238),
	   .D (n1183),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0194 (
	   .Q (_net_6135),
	   .D (n1178),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0193 (
	   .Q (net_7523),
	   .D (n1173),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0192 (
	   .Q (net_363),
	   .D (n1168),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0191 (
	   .Q (net_7611),
	   .D (n1163),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0190 (
	   .Q (net_6242),
	   .D (n1158),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0189 (
	   .Q (_net_6167),
	   .D (n1153),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0188 (
	   .Q (net_6677),
	   .D (n1148),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0187 (
	   .Q (net_6275),
	   .D (n1144),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0186 (
	   .Q (net_6986),
	   .D (n1140),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0185 (
	   .Q (_net_7299),
	   .D (n1135),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0184 (
	   .Q (net_6671),
	   .D (n1130),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0183 (
	   .Q (_net_7274),
	   .D (n1125),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0182 (
	   .Q (net_6847),
	   .D (n1121),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0181 (
	   .Q (net_6060),
	   .D (n1116),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0180 (
	   .Q (net_6379),
	   .D (n1111),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0179 (
	   .Q (_net_7412),
	   .D (n1106),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0178 (
	   .Q (net_6856),
	   .D (n1102),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0177 (
	   .Q (net_6901),
	   .D (n1097),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0176 (
	   .Q (net_6977),
	   .D (n1093),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0175 (
	   .Q (net_6832),
	   .D (n1089),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0174 (
	   .Q (net_6461),
	   .D (n1085),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0173 (
	   .Q (net_7010),
	   .D (n1081),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0172 (
	   .Q (net_7004),
	   .D (n1077),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0171 (
	   .Q (_net_6286),
	   .D (n1072),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0170 (
	   .Q (net_5992),
	   .D (n1067),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0169 (
	   .Q (net_6944),
	   .D (n1062),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0168 (
	   .Q (x657),
	   .D (n1058),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0167 (
	   .Q (net_351),
	   .D (n1053),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0166 (
	   .Q (_net_7578),
	   .D (n1049),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0165 (
	   .Q (_net_7281),
	   .D (n1044),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0164 (
	   .Q (_net_6220),
	   .D (n1039),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0163 (
	   .Q (net_7311),
	   .D (n1034),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0162 (
	   .Q (net_7334),
	   .D (n1029),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0161 (
	   .Q (_net_7447),
	   .D (n1024),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0160 (
	   .Q (net_6998),
	   .D (n1020),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0159 (
	   .Q (_net_6120),
	   .D (n1015),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0158 (
	   .Q (_net_7621),
	   .D (n1010),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0157 (
	   .Q (net_6392),
	   .D (n1005),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0156 (
	   .Q (net_391),
	   .D (n1000),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0155 (
	   .Q (_net_5856),
	   .D (n995),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0154 (
	   .Q (_net_7653),
	   .D (n990),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0153 (
	   .Q (_net_282),
	   .D (n985),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0152 (
	   .Q (net_6999),
	   .D (n981),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0151 (
	   .Q (net_150),
	   .D (n976),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0150 (
	   .Q (_net_7296),
	   .D (n971),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0149 (
	   .Q (net_204),
	   .D (n966),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0148 (
	   .Q (_net_7629),
	   .D (n961),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0147 (
	   .Q (net_7058),
	   .D (n956),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0146 (
	   .Q (net_6989),
	   .D (n953),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0145 (
	   .Q (_net_7809),
	   .D (n948),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0144 (
	   .Q (_net_5851),
	   .D (n944),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0143 (
	   .Q (net_6979),
	   .D (n940),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0142 (
	   .Q (net_7066),
	   .D (n935),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0141 (
	   .Q (_net_7632),
	   .D (n930),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0140 (
	   .Q (_net_7354),
	   .D (n925),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0139 (
	   .Q (net_6356),
	   .D (n920),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0138 (
	   .Q (net_6746),
	   .D (n916),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0137 (
	   .Q (net_7073),
	   .D (n911),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0136 (
	   .Q (net_7067),
	   .D (n907),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0135 (
	   .Q (_net_7439),
	   .D (n903),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0134 (
	   .Q (net_6739),
	   .D (n899),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0133 (
	   .Q (net_347),
	   .D (n894),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0132 (
	   .Q (net_6616),
	   .D (n890),
	   .CK (ck_net_4_12_a_2) );
   DFF_X1 l0131 (
	   .Q (_net_6008),
	   .D (n885),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0130 (
	   .Q (net_6646),
	   .D (n880),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0129 (
	   .Q (net_7312),
	   .D (n875),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0128 (
	   .Q (net_6815),
	   .D (n870),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0127 (
	   .Q (net_6711),
	   .D (n867),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0126 (
	   .Q (_net_6086),
	   .D (n862),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0125 (
	   .Q (net_6521),
	   .D (n857),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0124 (
	   .Q (net_7390),
	   .D (n854),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0123 (
	   .Q (net_171),
	   .D (n849),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0122 (
	   .Q (net_326),
	   .D (n844),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0121 (
	   .Q (net_6545),
	   .D (n839),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0120 (
	   .Q (net_220),
	   .D (n834),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0119 (
	   .Q (net_7396),
	   .D (n830),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0118 (
	   .Q (_net_120),
	   .D (n825),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0117 (
	   .Q (_net_121),
	   .D (n820),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0116 (
	   .Q (net_6260),
	   .D (n815),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0115 (
	   .Q (net_6400),
	   .D (n811),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0114 (
	   .Q (_net_7786),
	   .D (n806),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0113 (
	   .Q (net_7133),
	   .D (n802),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0112 (
	   .Q (net_7134),
	   .D (n798),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0111 (
	   .Q (net_7607),
	   .D (n793),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0110 (
	   .Q (_net_6012),
	   .D (n788),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0109 (
	   .Q (net_139),
	   .D (n783),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0108 (
	   .Q (net_6386),
	   .D (n779),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0107 (
	   .Q (net_6380),
	   .D (n774),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0106 (
	   .Q (_net_7732),
	   .D (n770),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0105 (
	   .Q (_net_113),
	   .D (n765),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0104 (
	   .Q (net_6468),
	   .D (n761),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0103 (
	   .Q (_net_6147),
	   .D (n756),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0102 (
	   .Q (net_7758),
	   .D (n751),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0101 (
	   .Q (net_235),
	   .D (n746),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0100 (
	   .Q (net_6213),
	   .D (n741),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0099 (
	   .Q (_net_6037),
	   .D (n736),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0098 (
	   .Q (x561),
	   .D (n732),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0097 (
	   .Q (net_236),
	   .D (n727),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0096 (
	   .Q (net_361),
	   .D (n722),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0095 (
	   .Q (net_7637),
	   .D (n718),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0094 (
	   .Q (net_7774),
	   .D (n713),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0093 (
	   .Q (_net_7300),
	   .D (n708),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0092 (
	   .Q (net_6323),
	   .D (n703),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0091 (
	   .Q (net_7645),
	   .D (n698),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0090 (
	   .Q (_net_7271),
	   .D (n693),
	   .CK (ck_net_4_9_b_1) );
   DFF_X1 l0089 (
	   .Q (_net_7330),
	   .D (n688),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0088 (
	   .Q (net_6491),
	   .D (n683),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0087 (
	   .Q (net_6653),
	   .D (n678),
	   .CK (ck_net_4_12_b_1) );
   DFF_X1 l0086 (
	   .Q (_net_6208),
	   .D (n673),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0085 (
	   .Q (net_6440),
	   .D (n669),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0084 (
	   .Q (net_6384),
	   .D (n664),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0083 (
	   .Q (net_160),
	   .D (n659),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0082 (
	   .Q (_net_7753),
	   .D (n654),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0081 (
	   .Q (_net_212),
	   .D (n649),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0080 (
	   .Q (_net_7094),
	   .D (n644),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0079 (
	   .Q (_net_7694),
	   .D (n639),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0078 (
	   .Q (net_7487),
	   .D (n634),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0077 (
	   .Q (_net_7441),
	   .D (n629),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0076 (
	   .Q (net_7246),
	   .D (n625),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0075 (
	   .Q (_net_6004),
	   .D (n620),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0074 (
	   .Q (net_7604),
	   .D (n615),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0073 (
	   .Q (net_6900),
	   .D (n610),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0072 (
	   .Q (_net_6210),
	   .D (n605),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0071 (
	   .Q (_net_7285),
	   .D (n600),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0070 (
	   .Q (net_7492),
	   .D (n595),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0069 (
	   .Q (net_365),
	   .D (n590),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0068 (
	   .Q (net_6373),
	   .D (n585),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0067 (
	   .Q (_net_7794),
	   .D (n580),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0066 (
	   .Q (net_7342),
	   .D (n576),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0065 (
	   .Q (net_6218),
	   .D (n571),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0064 (
	   .Q (net_6773),
	   .D (n566),
	   .CK (ck_net_4_18_b_1) );
   DFF_X1 l0063 (
	   .Q (_net_6294),
	   .D (n561),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0062 (
	   .Q (net_6791),
	   .D (n556),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0061 (
	   .Q (x14),
	   .D (n553),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0060 (
	   .Q (_net_5965),
	   .D (n548),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0059 (
	   .Q (_net_7316),
	   .D (n543),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0058 (
	   .Q (_net_7603),
	   .D (n538),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0057 (
	   .Q (_net_6104),
	   .D (n533),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0056 (
	   .Q (_net_7689),
	   .D (n528),
	   .CK (ck_net_4_17_a_1) );
   DFF_X1 l0055 (
	   .Q (_net_6079),
	   .D (n523),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0054 (
	   .Q (net_7369),
	   .D (n518),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0053 (
	   .Q (net_6691),
	   .D (n513),
	   .CK (ck_net_4_14_a_2) );
   DFF_X1 l0052 (
	   .Q (net_6308),
	   .D (n508),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0051 (
	   .Q (net_6267),
	   .D (n503),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0050 (
	   .Q (_net_6194),
	   .D (n498),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0049 (
	   .Q (net_7224),
	   .D (n493),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0048 (
	   .Q (net_7196),
	   .D (n488),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0047 (
	   .Q (net_6870),
	   .D (n484),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0046 (
	   .Q (net_6783),
	   .D (n479),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0045 (
	   .Q (net_362),
	   .D (n474),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0044 (
	   .Q (net_7388),
	   .D (n470),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0043 (
	   .Q (_net_6100),
	   .D (n465),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0042 (
	   .Q (_net_7355),
	   .D (n460),
	   .CK (ck_net_4_8_b_1) );
   DFF_X1 l0041 (
	   .Q (net_6628),
	   .D (n455),
	   .CK (ck_net_4_13_b_1) );
   DFF_X1 l0040 (
	   .Q (net_7802),
	   .D (n451),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0039 (
	   .Q (_net_6150),
	   .D (n447),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0038 (
	   .Q (net_7000),
	   .D (n443),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0037 (
	   .Q (net_6510),
	   .D (n438),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0036 (
	   .Q (net_7713),
	   .D (n434),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0035 (
	   .Q (net_6803),
	   .D (n429),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0034 (
	   .Q (net_6514),
	   .D (n424),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0033 (
	   .Q (net_7525),
	   .D (n420),
	   .CK (ck_net_4_16_a_1) );
   DFF_X1 l0032 (
	   .Q (net_7062),
	   .D (n415),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0031 (
	   .Q (net_6313),
	   .D (n410),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0030 (
	   .Q (net_6396),
	   .D (n405),
	   .CK (ck_net_4_10_b_1) );
   DFF_X1 l0029 (
	   .Q (_net_7595),
	   .D (n400),
	   .CK (ck_net_4_15_a_2) );
   DFF_X1 l0028 (
	   .Q (net_7055),
	   .D (n395),
	   .CK (ck_net_4_11_b_1) );
   DFF_X1 l0027 (
	   .Q (_net_6088),
	   .D (n390),
	   .CK (ck_net_4_14_b_1) );
   DFF_X1 l0026 (
	   .Q (_net_6404),
	   .D (n385),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0025 (
	   .Q (_net_298),
	   .D (n380),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0024 (
	   .Q (_net_7252),
	   .D (n375),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0023 (
	   .Q (_net_7474),
	   .D (n370),
	   .CK (ck_net_4_18_a_1) );
   DFF_X1 l0022 (
	   .Q (net_6996),
	   .D (n366),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0021 (
	   .Q (net_6784),
	   .D (n361),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0020 (
	   .Q (net_7114),
	   .D (n357),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0019 (
	   .Q (_net_7800),
	   .D (n352),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0018 (
	   .Q (net_6474),
	   .D (n349),
	   .CK (ck_net_4_19_a_2) );
   DFF_X1 l0017 (
	   .Q (net_6256),
	   .D (n344),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0016 (
	   .Q (net_6364),
	   .D (n339),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0015 (
	   .Q (net_6227),
	   .D (n334),
	   .CK (ck_net_4_7_a_1) );
   DFF_X1 l0014 (
	   .Q (_net_6062),
	   .D (n329),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0013 (
	   .Q (net_7204),
	   .D (n324),
	   .CK (ck_net_4_22_b_1) );
   DFF_X1 l0012 (
	   .Q (_net_175),
	   .D (n319),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0011 (
	   .Q (_net_7481),
	   .D (n314),
	   .CK (ck_net_4_16_b_1) );
   DFF_X1 l0010 (
	   .Q (net_6704),
	   .D (n310),
	   .CK (ck_net_4_17_b_1) );
   DFF_X1 l0009 (
	   .Q (net_7222),
	   .D (n305),
	   .CK (ck_net_4_21_b_1) );
   DFF_X1 l0008 (
	   .Q (_net_6133),
	   .D (n300),
	   .CK (ck_net_4_7_b_1) );
   DFF_X1 l0007 (
	   .Q (_net_6032),
	   .D (n295),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0006 (
	   .Q (net_6453),
	   .D (n291),
	   .CK (ck_net_4_20_b_1) );
   DFF_X1 l0005 (
	   .Q (net_6300),
	   .D (n286),
	   .CK (ck_net_1_0_b_2) );
   DFF_X1 l0004 (
	   .Q (_net_6082),
	   .D (n281),
	   .CK (ck_net_4_19_b_1) );
   DFF_X1 l0003 (
	   .Q (net_6907),
	   .D (n276),
	   .CK (ck_net_1_0_a_2) );
   DFF_X1 l0002 (
	   .Q (net_254),
	   .D (n271),
	   .CK (ck_net_4_15_b_1) );
   DFF_X1 l0001 (
	   .Q (net_249),
	   .D (n266),
	   .CK (ck_net_4_15_b_1) );
   CLKBUF_X1 g5608 (
	   .Z (n10158),
	   .A (_net_7806) );
   CLKBUF_X1 g5607 (
	   .Z (n10154),
	   .A (net_7807) );
   OAI21_X1 g5606 (
	   .ZN (n10150),
	   .B2 (new_n7692_),
	   .B1 (new_n11683_),
	   .A (new_n12336_) );
   NAND2_X1 g5605 (
	   .ZN (new_n12336_),
	   .A2 (new_n7690_),
	   .A1 (new_n8034_) );
   NOR2_X1 g5604 (
	   .ZN (n10145),
	   .A2 (new_n7602_),
	   .A1 (new_n8675_) );
   CLKBUF_X1 g5603 (
	   .Z (n10141),
	   .A (x1595) );
   NAND3_X1 g5602 (
	   .ZN (n10137),
	   .A3 (new_n12332_),
	   .A2 (new_n12331_),
	   .A1 (new_n12327_) );
   AOI22_X1 g5601 (
	   .ZN (new_n12332_),
	   .B2 (net_7219),
	   .B1 (new_n7844_),
	   .A2 (new_n9781_),
	   .A1 (new_n7837_) );
   AND3_X1 g5600 (
	   .ZN (new_n12331_),
	   .A3 (new_n12330_),
	   .A2 (new_n12329_),
	   .A1 (new_n12328_) );
   NAND2_X1 g5599 (
	   .ZN (new_n12330_),
	   .A2 (_net_6176),
	   .A1 (new_n7693_) );
   NAND2_X1 g5598 (
	   .ZN (new_n12329_),
	   .A2 (new_n7700_1_),
	   .A1 (new_n11639_) );
   NAND2_X1 g5597 (
	   .ZN (new_n12328_),
	   .A2 (new_n7689_),
	   .A1 (new_n8060_) );
   AND3_X1 g5596 (
	   .ZN (new_n12327_),
	   .A3 (new_n12326_),
	   .A2 (new_n12325_),
	   .A1 (new_n12324_) );
   NAND4_X1 g5595 (
	   .ZN (new_n12326_),
	   .A4 (new_n7678_),
	   .A3 (net_7187),
	   .A2 (_net_7227),
	   .A1 (new_n7812_) );
   NAND4_X1 g5594 (
	   .ZN (new_n12325_),
	   .A4 (new_n7683_),
	   .A3 (net_7123),
	   .A2 (_net_7227),
	   .A1 (new_n7816_) );
   NAND4_X1 g5593 (
	   .ZN (new_n12324_),
	   .A4 (new_n7681_1_),
	   .A3 (net_7155),
	   .A2 (_net_7227),
	   .A1 (new_n7813_) );
   CLKBUF_X1 g5592 (
	   .Z (n10132),
	   .A (_net_7805) );
   OAI21_X1 g5591 (
	   .ZN (n10128),
	   .B2 (new_n7101_),
	   .B1 (new_n11663_),
	   .A (new_n12321_) );
   NAND2_X1 g5590 (
	   .ZN (new_n12321_),
	   .A2 (new_n10131_),
	   .A1 (new_n7100_) );
   CLKBUF_X1 g5589 (
	   .Z (n10124),
	   .A (_net_7811) );
   CLKBUF_X1 g5588 (
	   .Z (n10120),
	   .A (_net_7815) );
   NAND2_X1 g5587 (
	   .ZN (n10116),
	   .A2 (new_n12317_),
	   .A1 (new_n12316_) );
   AOI22_X1 g5586 (
	   .ZN (new_n12317_),
	   .B2 (new_n6751_),
	   .B1 (_net_7570),
	   .A2 (_net_7666),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g5585 (
	   .ZN (new_n12316_),
	   .B2 (_net_7602),
	   .B1 (new_n7350_),
	   .A2 (new_n6746_1_),
	   .A1 (_net_7634) );
   CLKBUF_X1 g5584 (
	   .Z (n10112),
	   .A (net_7112) );
   CLKBUF_X1 g5583 (
	   .Z (n10107),
	   .A (_net_7818) );
   CLKBUF_X1 g5582 (
	   .Z (n10103),
	   .A (_net_7815) );
   OAI21_X1 g5581 (
	   .ZN (n10099),
	   .B2 (new_n6897_),
	   .B1 (new_n8696_),
	   .A (new_n12311_) );
   NAND2_X1 g5580 (
	   .ZN (new_n12311_),
	   .A2 (new_n7595_),
	   .A1 (new_n6896_) );
   OAI21_X1 g5579 (
	   .ZN (n10094),
	   .B2 (new_n6949_),
	   .B1 (new_n12309_),
	   .A (new_n12308_) );
   INV_X1 g5578 (
	   .ZN (new_n12309_),
	   .A (_net_7264) );
   NAND2_X1 g5577 (
	   .ZN (new_n12308_),
	   .A2 (new_n7531_),
	   .A1 (new_n6948_) );
   NAND3_X1 g5576 (
	   .ZN (n10089),
	   .A3 (new_n12306_),
	   .A2 (new_n12305_),
	   .A1 (new_n12301_) );
   AOI22_X1 g5575 (
	   .ZN (new_n12306_),
	   .B2 (net_7226),
	   .B1 (new_n7844_),
	   .A2 (new_n10495_),
	   .A1 (new_n7837_) );
   AND3_X1 g5574 (
	   .ZN (new_n12305_),
	   .A3 (new_n12304_),
	   .A2 (new_n12303_),
	   .A1 (new_n12302_) );
   NAND2_X1 g5573 (
	   .ZN (new_n12304_),
	   .A2 (_net_6183),
	   .A1 (new_n7693_) );
   NAND2_X1 g5572 (
	   .ZN (new_n12303_),
	   .A2 (new_n7689_),
	   .A1 (new_n9109_) );
   NAND2_X1 g5571 (
	   .ZN (new_n12302_),
	   .A2 (new_n7701_),
	   .A1 (new_n8553_) );
   AND3_X1 g5570 (
	   .ZN (new_n12301_),
	   .A3 (new_n12300_),
	   .A2 (new_n12299_),
	   .A1 (new_n12298_) );
   NAND4_X1 g5569 (
	   .ZN (new_n12300_),
	   .A4 (new_n7678_),
	   .A3 (_net_7227),
	   .A2 (net_7194),
	   .A1 (new_n7812_) );
   NAND4_X1 g5568 (
	   .ZN (new_n12299_),
	   .A4 (new_n7683_),
	   .A3 (net_7130),
	   .A2 (_net_7227),
	   .A1 (new_n7816_) );
   NAND4_X1 g5567 (
	   .ZN (new_n12298_),
	   .A4 (new_n7681_1_),
	   .A3 (net_7162),
	   .A2 (_net_7227),
	   .A1 (new_n7813_) );
   NAND4_X1 g5566 (
	   .ZN (n10084),
	   .A4 (new_n12296_),
	   .A3 (new_n12295_),
	   .A2 (new_n12294_),
	   .A1 (new_n12293_) );
   AOI22_X1 g5565 (
	   .ZN (new_n12296_),
	   .B2 (_net_6131),
	   .B1 (new_n6869_),
	   .A2 (new_n6854_),
	   .A1 (new_n6860_1_) );
   NAND2_X1 g5564 (
	   .ZN (new_n12295_),
	   .A2 (new_n12127_),
	   .A1 (new_n9255_) );
   NAND2_X1 g5563 (
	   .ZN (new_n12294_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n6876_1_) );
   NAND2_X1 g5562 (
	   .ZN (new_n12293_),
	   .A2 (new_n6879_),
	   .A1 (new_n10783_) );
   OAI211_X1 g5561 (
	   .ZN (n10079),
	   .C2 (new_n12291_),
	   .C1 (new_n7858_1_),
	   .B (new_n12290_),
	   .A (new_n12289_) );
   INV_X1 g5560 (
	   .ZN (new_n12291_),
	   .A (new_n8908_1_) );
   NAND2_X1 g5559 (
	   .ZN (new_n12290_),
	   .A2 (_net_6555),
	   .A1 (new_n6813_1_) );
   OAI21_X1 g5558 (
	   .ZN (new_n12289_),
	   .B2 (new_n7861_),
	   .B1 (new_n7860_),
	   .A (new_n6764_) );
   OAI21_X1 g5557 (
	   .ZN (n10074),
	   .B2 (new_n6949_),
	   .B1 (new_n12287_),
	   .A (new_n12286_) );
   INV_X1 g5556 (
	   .ZN (new_n12287_),
	   .A (_net_7251) );
   NAND2_X1 g5555 (
	   .ZN (new_n12286_),
	   .A2 (new_n7773_1_),
	   .A1 (new_n6948_) );
   CLKBUF_X1 g5554 (
	   .Z (n10070),
	   .A (net_6884) );
   NAND3_X1 g5553 (
	   .ZN (n10066),
	   .A3 (new_n12283_),
	   .A2 (new_n12282_),
	   .A1 (new_n12274_) );
   OR2_X1 g5552 (
	   .ZN (new_n12283_),
	   .A2 (new_n7508_),
	   .A1 (new_n7362_) );
   NOR3_X1 g5551 (
	   .ZN (new_n12282_),
	   .A3 (new_n12281_),
	   .A2 (new_n12277_),
	   .A1 (new_n12275_) );
   NAND3_X1 g5550 (
	   .ZN (new_n12281_),
	   .A3 (new_n12280_),
	   .A2 (new_n12279_),
	   .A1 (new_n12278_) );
   NAND4_X1 g5549 (
	   .ZN (new_n12280_),
	   .A4 (net_164),
	   .A3 (x1231),
	   .A2 (new_n7394_),
	   .A1 (new_n7392_) );
   NAND3_X1 g5548 (
	   .ZN (new_n12279_),
	   .A3 (_net_201),
	   .A2 (new_n7388_),
	   .A1 (new_n7386_1_) );
   NAND3_X1 g5547 (
	   .ZN (new_n12278_),
	   .A3 (net_238),
	   .A2 (new_n7382_),
	   .A1 (new_n7380_) );
   OAI22_X1 g5546 (
	   .ZN (new_n12277_),
	   .B2 (new_n7377_),
	   .B1 (new_n9371_),
	   .A2 (new_n12276_),
	   .A1 (new_n7374_) );
   INV_X1 g5545 (
	   .ZN (new_n12276_),
	   .A (_net_122) );
   AND4_X1 g5544 (
	   .ZN (new_n12275_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7357_),
	   .A1 (_net_6039) );
   NOR2_X1 g5543 (
	   .ZN (new_n12274_),
	   .A2 (new_n12273_),
	   .A1 (new_n12272_) );
   NOR2_X1 g5542 (
	   .ZN (new_n12273_),
	   .A2 (new_n6983_),
	   .A1 (new_n7365_) );
   NOR2_X1 g5541 (
	   .ZN (new_n12272_),
	   .A2 (new_n12271_),
	   .A1 (new_n9215_1_) );
   INV_X1 g5540 (
	   .ZN (new_n12271_),
	   .A (_net_7699) );
   NOR2_X1 g5539 (
	   .ZN (n10061),
	   .A2 (x1034),
	   .A1 (new_n12269_) );
   NAND2_X1 g5538 (
	   .ZN (new_n12269_),
	   .A2 (_net_6001),
	   .A1 (n6643) );
   AND2_X1 g5537 (
	   .ZN (n10056),
	   .A2 (net_383),
	   .A1 (new_n7262_) );
   OAI21_X1 g5536 (
	   .ZN (n10052),
	   .B2 (new_n7252_1_),
	   .B1 (new_n11047_),
	   .A (new_n12266_) );
   NAND2_X1 g5535 (
	   .ZN (new_n12266_),
	   .A2 (new_n8133_),
	   .A1 (new_n7251_) );
   CLKBUF_X1 g5534 (
	   .Z (n10047),
	   .A (_net_6155) );
   AND2_X1 g5533 (
	   .ZN (n10042),
	   .A2 (_net_6202),
	   .A1 (new_n7235_1_) );
   MUX2_X1 g5532 (
	   .Z (n10037),
	   .S (new_n7436_),
	   .B (_net_6017),
	   .A (_net_7817) );
   MUX2_X1 g5531 (
	   .Z (n10032),
	   .S (new_n10364_),
	   .B (_net_7582),
	   .A (n3604) );
   CLKBUF_X1 g5530 (
	   .Z (n10028),
	   .A (net_6879) );
   CLKBUF_X1 g5529 (
	   .Z (n10023),
	   .A (net_130) );
   MUX2_X1 g5528 (
	   .Z (n10019),
	   .S (new_n7537_),
	   .B (_net_267),
	   .A (_net_7793) );
   CLKBUF_X1 g5527 (
	   .Z (n10014),
	   .A (x1351) );
   CLKBUF_X1 g5526 (
	   .Z (n10010),
	   .A (net_7802) );
   CLKBUF_X1 g5525 (
	   .Z (n10006),
	   .A (_net_6062) );
   CLKBUF_X1 g5524 (
	   .Z (n10001),
	   .A (_net_7812) );
   MUX2_X1 g5523 (
	   .Z (n9997),
	   .S (new_n7284_1_),
	   .B (_net_7717),
	   .A (_net_7819) );
   CLKBUF_X1 g5522 (
	   .Z (n9992),
	   .A (_net_7805) );
   CLKBUF_X1 g5521 (
	   .Z (n9988),
	   .A (_net_7805) );
   CLKBUF_X1 g5520 (
	   .Z (n9985),
	   .A (net_6380) );
   NOR3_X1 g5519 (
	   .ZN (n9981),
	   .A3 (new_n12249_),
	   .A2 (new_n10598_),
	   .A1 (new_n7449_) );
   NOR2_X1 g5518 (
	   .ZN (new_n12249_),
	   .A2 (_net_7788),
	   .A1 (new_n10597_) );
   CLKBUF_X1 g5517 (
	   .Z (n9976),
	   .A (net_6057) );
   NAND3_X1 g5516 (
	   .ZN (n9971),
	   .A3 (new_n12246_),
	   .A2 (new_n12242_),
	   .A1 (new_n12241_) );
   AND3_X1 g5515 (
	   .ZN (new_n12246_),
	   .A3 (new_n12245_),
	   .A2 (new_n12244_),
	   .A1 (new_n12243_) );
   NAND2_X1 g5514 (
	   .ZN (new_n12245_),
	   .A2 (_net_6076),
	   .A1 (new_n6812_) );
   NAND2_X1 g5513 (
	   .ZN (new_n12244_),
	   .A2 (new_n6800_),
	   .A1 (new_n9275_) );
   NAND2_X1 g5512 (
	   .ZN (new_n12243_),
	   .A2 (new_n6809_1_),
	   .A1 (new_n9282_1_) );
   AOI22_X1 g5511 (
	   .ZN (new_n12242_),
	   .B2 (new_n10625_),
	   .B1 (new_n6783_1_),
	   .A2 (new_n6779_1_),
	   .A1 (net_6544) );
   AND3_X1 g5510 (
	   .ZN (new_n12241_),
	   .A3 (new_n12240_),
	   .A2 (new_n12239_),
	   .A1 (new_n12238_) );
   NAND4_X1 g5509 (
	   .ZN (new_n12240_),
	   .A4 (new_n6775_),
	   .A3 (_net_6552),
	   .A2 (net_6512),
	   .A1 (new_n6763_) );
   NAND4_X1 g5508 (
	   .ZN (new_n12239_),
	   .A4 (new_n6770_1_),
	   .A3 (_net_6552),
	   .A2 (net_6448),
	   .A1 (new_n6772_) );
   NAND4_X1 g5507 (
	   .ZN (new_n12238_),
	   .A4 (new_n6767_),
	   .A3 (_net_6552),
	   .A2 (net_6480),
	   .A1 (new_n6764_) );
   OAI21_X1 g5506 (
	   .ZN (n9966),
	   .B2 (new_n7646_),
	   .B1 (new_n12236_),
	   .A (new_n12235_) );
   INV_X1 g5505 (
	   .ZN (new_n12236_),
	   .A (_net_7402) );
   NAND2_X1 g5504 (
	   .ZN (new_n12235_),
	   .A2 (new_n7991_),
	   .A1 (new_n7645_) );
   CLKBUF_X1 g5503 (
	   .Z (n9961),
	   .A (_net_7804) );
   CLKBUF_X1 g5502 (
	   .Z (n9957),
	   .A (net_6389) );
   NAND2_X1 g5501 (
	   .ZN (n9953),
	   .A2 (n4304),
	   .A1 (new_n7422_1_) );
   OAI21_X1 g5500 (
	   .ZN (n9949),
	   .B2 (new_n7101_),
	   .B1 (new_n11406_),
	   .A (new_n12230_) );
   NAND2_X1 g5499 (
	   .ZN (new_n12230_),
	   .A2 (new_n6954_),
	   .A1 (new_n7100_) );
   CLKBUF_X1 g5498 (
	   .Z (n9944),
	   .A (_net_6174) );
   OAI21_X1 g5497 (
	   .ZN (n9939),
	   .B2 (new_n12227_),
	   .B1 (new_n7950_1_),
	   .A (new_n11987_) );
   INV_X1 g5496 (
	   .ZN (new_n12227_),
	   .A (_net_226) );
   CLKBUF_X1 g5495 (
	   .Z (n9935),
	   .A (net_6465) );
   CLKBUF_X1 g5494 (
	   .Z (n9930),
	   .A (net_6393) );
   CLKBUF_X1 g5493 (
	   .Z (n9926),
	   .A (net_6389) );
   CLKBUF_X1 g5492 (
	   .Z (n9923),
	   .A (net_6719) );
   CLKBUF_X1 g5491 (
	   .Z (n9918),
	   .A (x1580) );
   CLKBUF_X1 g5490 (
	   .Z (n9914),
	   .A (_net_7819) );
   CLKBUF_X1 g5489 (
	   .Z (n9911),
	   .A (net_6446) );
   NAND4_X1 g5488 (
	   .ZN (n9907),
	   .A4 (new_n12218_),
	   .A3 (new_n12217_),
	   .A2 (new_n12216_),
	   .A1 (new_n12215_) );
   NAND4_X1 g5487 (
	   .ZN (new_n12218_),
	   .A4 (net_7711),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7399_) );
   NAND4_X1 g5486 (
	   .ZN (new_n12217_),
	   .A4 (new_n7364_),
	   .A3 (_net_6010),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   NAND4_X1 g5485 (
	   .ZN (new_n12216_),
	   .A4 (_net_293),
	   .A3 (x1286),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR2_X1 g5484 (
	   .ZN (new_n12215_),
	   .A2 (new_n12214_),
	   .A1 (new_n12213_) );
   AND2_X1 g5483 (
	   .ZN (new_n12214_),
	   .A2 (net_7740),
	   .A1 (new_n7934_) );
   NAND4_X1 g5482 (
	   .ZN (new_n12213_),
	   .A4 (new_n12212_),
	   .A3 (new_n12211_),
	   .A2 (new_n12210_),
	   .A1 (new_n12209_) );
   NAND4_X1 g5481 (
	   .ZN (new_n12212_),
	   .A4 (_net_176),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g5480 (
	   .ZN (new_n12211_),
	   .A3 (_net_213),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g5479 (
	   .ZN (new_n12210_),
	   .A3 (net_250),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   NAND4_X1 g5478 (
	   .ZN (new_n12209_),
	   .A4 (new_n7354_1_),
	   .A3 (net_150),
	   .A2 (x1261),
	   .A1 (new_n7370_) );
   CLKBUF_X1 g5477 (
	   .Z (n9902),
	   .A (_net_7798) );
   CLKBUF_X1 g5476 (
	   .Z (n9899),
	   .A (net_6752) );
   OAI21_X1 g5475 (
	   .ZN (n9894),
	   .B2 (new_n12205_),
	   .B1 (new_n10359_),
	   .A (new_n12204_) );
   INV_X1 g5474 (
	   .ZN (new_n12205_),
	   .A (_net_225) );
   INV_X1 g5473 (
	   .ZN (new_n12204_),
	   .A (_net_287) );
   NAND4_X1 g5472 (
	   .ZN (n9889),
	   .A4 (new_n12202_),
	   .A3 (new_n12201_),
	   .A2 (new_n12200_),
	   .A1 (new_n12199_) );
   AOI22_X1 g5471 (
	   .ZN (new_n12202_),
	   .B2 (_net_6111),
	   .B1 (new_n7210_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n10836_) );
   NAND2_X1 g5470 (
	   .ZN (new_n12201_),
	   .A2 (new_n7587_),
	   .A1 (new_n10824_) );
   NAND2_X1 g5469 (
	   .ZN (new_n12200_),
	   .A2 (new_n11561_),
	   .A1 (new_n7556_) );
   NAND2_X1 g5468 (
	   .ZN (new_n12199_),
	   .A2 (new_n7565_),
	   .A1 (new_n8271_1_) );
   CLKBUF_X1 g5467 (
	   .Z (n9885),
	   .A (net_7109) );
   OAI22_X1 g5466 (
	   .ZN (n9880),
	   .B2 (new_n9435_),
	   .B1 (new_n10159_),
	   .A2 (new_n12196_),
	   .A1 (new_n12195_) );
   XNOR2_X1 g5465 (
	   .ZN (new_n12196_),
	   .B (new_n9435_),
	   .A (new_n9675_) );
   INV_X1 g5464 (
	   .ZN (new_n12195_),
	   .A (new_n9673_1_) );
   CLKBUF_X1 g5463 (
	   .Z (n9875),
	   .A (_net_7806) );
   CLKBUF_X1 g5462 (
	   .Z (n9871),
	   .A (_net_7797) );
   CLKBUF_X1 g5461 (
	   .Z (n9867),
	   .A (_net_7811) );
   NOR3_X1 g5460 (
	   .ZN (n9863),
	   .A3 (new_n12190_),
	   .A2 (new_n7090_),
	   .A1 (new_n10641_) );
   AOI21_X1 g5459 (
	   .ZN (new_n12190_),
	   .B2 (_net_5979),
	   .B1 (net_7096),
	   .A (_net_7097) );
   OAI21_X1 g5458 (
	   .ZN (n9858),
	   .B2 (new_n9305_),
	   .B1 (new_n12188_),
	   .A (new_n6963_) );
   NOR2_X1 g5457 (
	   .ZN (new_n12188_),
	   .A2 (_net_6407),
	   .A1 (new_n9935_1_) );
   AND2_X1 g5456 (
	   .ZN (n9853),
	   .A2 (net_382),
	   .A1 (new_n7262_) );
   AOI21_X1 g5455 (
	   .ZN (n9849),
	   .B2 (new_n7739_),
	   .B1 (new_n12185_),
	   .A (new_n12184_) );
   INV_X1 g5454 (
	   .ZN (new_n12185_),
	   .A (_net_7421) );
   NOR2_X1 g5453 (
	   .ZN (new_n12184_),
	   .A2 (n1277),
	   .A1 (new_n7738_) );
   CLKBUF_X1 g5452 (
	   .Z (n9844),
	   .A (net_6387) );
   CLKBUF_X1 g5451 (
	   .Z (n9840),
	   .A (net_6396) );
   CLKBUF_X1 g5450 (
	   .Z (n9837),
	   .A (net_7122) );
   CLKBUF_X1 g5449 (
	   .Z (n9833),
	   .A (net_7135) );
   AND2_X1 g5448 (
	   .ZN (n9828),
	   .A2 (net_380),
	   .A1 (new_n7262_) );
   OAI211_X1 g5447 (
	   .ZN (n9824),
	   .C2 (new_n12177_),
	   .C1 (new_n11207_),
	   .B (new_n12176_),
	   .A (new_n12175_) );
   NOR2_X1 g5446 (
	   .ZN (new_n12177_),
	   .A2 (new_n7249_1_),
	   .A1 (new_n7219_) );
   NAND3_X1 g5445 (
	   .ZN (new_n12176_),
	   .A3 (_net_267),
	   .A2 (_net_7383),
	   .A1 (new_n9619_) );
   NAND4_X1 g5444 (
	   .ZN (new_n12175_),
	   .A4 (new_n12174_),
	   .A3 (new_n12164_),
	   .A2 (new_n7102_1_),
	   .A1 (new_n11205_) );
   OAI21_X1 g5443 (
	   .ZN (new_n12174_),
	   .B2 (new_n6943_1_),
	   .B1 (new_n7248_),
	   .A (new_n7218_) );
   AOI21_X1 g5442 (
	   .ZN (n9819),
	   .B2 (new_n6892_),
	   .B1 (_net_7533),
	   .A (new_n12172_) );
   OAI21_X1 g5441 (
	   .ZN (new_n12172_),
	   .B2 (_net_7533),
	   .B1 (new_n6892_),
	   .A (_net_278) );
   NOR2_X1 g5440 (
	   .ZN (n9814),
	   .A2 (x1062),
	   .A1 (new_n12170_) );
   AOI21_X1 g5439 (
	   .ZN (new_n12170_),
	   .B2 (net_7772),
	   .B1 (new_n11512_),
	   .A (_net_5859) );
   CLKBUF_X1 g5438 (
	   .Z (n9809),
	   .A (net_6388) );
   CLKBUF_X1 g5437 (
	   .Z (n9805),
	   .A (net_6399) );
   AOI221_X4 g5436 (
	   .ZN (n9801),
	   .C2 (new_n12163_),
	   .C1 (new_n12166_),
	   .B2 (new_n6941_),
	   .B1 (new_n12165_),
	   .A (new_n8193_) );
   NAND2_X1 g5435 (
	   .ZN (new_n12166_),
	   .A2 (new_n7098_1_),
	   .A1 (new_n6945_) );
   OAI21_X1 g5434 (
	   .ZN (new_n12165_),
	   .B2 (new_n12164_),
	   .B1 (new_n12163_),
	   .A (new_n12162_) );
   NAND3_X1 g5433 (
	   .ZN (new_n12164_),
	   .A3 (_net_7383),
	   .A2 (_net_7381),
	   .A1 (_net_7382) );
   INV_X1 g5432 (
	   .ZN (new_n12163_),
	   .A (_net_7384) );
   NAND3_X1 g5431 (
	   .ZN (new_n12162_),
	   .A3 (_net_7384),
	   .A2 (new_n7098_1_),
	   .A1 (new_n6951_) );
   CLKBUF_X1 g5430 (
	   .Z (n9796),
	   .A (_net_7810) );
   MUX2_X1 g5429 (
	   .Z (n9792),
	   .S (new_n7436_),
	   .B (_net_5989),
	   .A (_net_7798) );
   MUX2_X1 g5428 (
	   .Z (n9787),
	   .S (new_n10364_),
	   .B (_net_7566),
	   .A (new_n9405_1_) );
   CLKBUF_X1 g5427 (
	   .Z (n9783),
	   .A (net_7027) );
   MUX2_X1 g5426 (
	   .Z (n9773),
	   .S (new_n7436_),
	   .B (_net_6002),
	   .A (_net_7808) );
   OAI21_X1 g5425 (
	   .ZN (n9768),
	   .B2 (new_n7252_1_),
	   .B1 (new_n10730_),
	   .A (new_n12155_) );
   NAND2_X1 g5424 (
	   .ZN (new_n12155_),
	   .A2 (new_n7773_1_),
	   .A1 (new_n7251_) );
   MUX2_X1 g5423 (
	   .Z (n9763),
	   .S (new_n10364_),
	   .B (_net_7576),
	   .A (n2404) );
   AND2_X1 g5422 (
	   .ZN (n9758),
	   .A2 (net_375),
	   .A1 (new_n7262_) );
   NOR2_X1 g5421 (
	   .ZN (n9754),
	   .A2 (new_n7648_),
	   .A1 (new_n7035_) );
   CLKBUF_X1 g5420 (
	   .Z (n9750),
	   .A (_net_7795) );
   CLKBUF_X1 g5419 (
	   .Z (n9746),
	   .A (_net_7812) );
   OAI221_X1 g5418 (
	   .ZN (n9742),
	   .C2 (new_n6920_),
	   .C1 (new_n10414_),
	   .B2 (new_n6917_),
	   .B1 (new_n7533_),
	   .A (new_n12148_) );
   AOI22_X1 g5417 (
	   .ZN (new_n12148_),
	   .B2 (_net_7264),
	   .B1 (new_n10556_),
	   .A2 (_net_7328),
	   .A1 (new_n10555_) );
   CLKBUF_X1 g5416 (
	   .Z (n9737),
	   .A (x1398) );
   XNOR2_X1 g5415 (
	   .ZN (n9733),
	   .B (new_n12145_),
	   .A (new_n9462_1_) );
   NAND2_X1 g5414 (
	   .ZN (new_n12145_),
	   .A2 (net_7378),
	   .A1 (new_n7248_) );
   CLKBUF_X1 g5413 (
	   .Z (n9729),
	   .A (net_6472) );
   CLKBUF_X1 g5412 (
	   .Z (n9724),
	   .A (_net_6162) );
   NAND3_X1 g5411 (
	   .ZN (n9719),
	   .A3 (new_n12141_),
	   .A2 (new_n12140_),
	   .A1 (new_n12136_) );
   AOI22_X1 g5410 (
	   .ZN (new_n12141_),
	   .B2 (net_7217),
	   .B1 (new_n7844_),
	   .A2 (new_n9787_1_),
	   .A1 (new_n7837_) );
   AND3_X1 g5409 (
	   .ZN (new_n12140_),
	   .A3 (new_n12139_),
	   .A2 (new_n12138_),
	   .A1 (new_n12137_) );
   NAND2_X1 g5408 (
	   .ZN (new_n12139_),
	   .A2 (_net_6174),
	   .A1 (new_n7693_) );
   NAND2_X1 g5407 (
	   .ZN (new_n12138_),
	   .A2 (new_n7700_1_),
	   .A1 (new_n9781_) );
   NAND2_X1 g5406 (
	   .ZN (new_n12137_),
	   .A2 (new_n7689_),
	   .A1 (new_n11639_) );
   AND3_X1 g5405 (
	   .ZN (new_n12136_),
	   .A3 (new_n12135_),
	   .A2 (new_n12134_),
	   .A1 (new_n12133_) );
   NAND4_X1 g5404 (
	   .ZN (new_n12135_),
	   .A4 (new_n7678_),
	   .A3 (_net_7227),
	   .A2 (net_7185),
	   .A1 (new_n7812_) );
   NAND4_X1 g5403 (
	   .ZN (new_n12134_),
	   .A4 (new_n7683_),
	   .A3 (_net_7227),
	   .A2 (net_7121),
	   .A1 (new_n7816_) );
   NAND4_X1 g5402 (
	   .ZN (new_n12133_),
	   .A4 (new_n7681_1_),
	   .A3 (_net_7227),
	   .A2 (net_7153),
	   .A1 (new_n7813_) );
   NAND3_X1 g5401 (
	   .ZN (n9714),
	   .A3 (new_n12131_),
	   .A2 (new_n12130_),
	   .A1 (new_n12121_) );
   AOI22_X1 g5400 (
	   .ZN (new_n12131_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6956),
	   .A2 (new_n8451_1_),
	   .A1 (new_n6879_) );
   AND3_X1 g5399 (
	   .ZN (new_n12130_),
	   .A3 (new_n12129_),
	   .A2 (new_n12128_),
	   .A1 (new_n12122_) );
   NAND2_X1 g5398 (
	   .ZN (new_n12129_),
	   .A2 (_net_6143),
	   .A1 (new_n6868_) );
   NAND2_X1 g5397 (
	   .ZN (new_n12128_),
	   .A2 (new_n6853_),
	   .A1 (new_n12127_) );
   NAND4_X1 g5396 (
	   .ZN (new_n12127_),
	   .A4 (new_n12126_),
	   .A3 (new_n12125_),
	   .A2 (new_n12124_),
	   .A1 (new_n12123_) );
   NAND3_X1 g5395 (
	   .ZN (new_n12126_),
	   .A3 (_net_6958),
	   .A2 (_net_6959),
	   .A1 (net_6944) );
   NAND3_X1 g5394 (
	   .ZN (new_n12125_),
	   .A3 (_net_6959),
	   .A2 (net_6912),
	   .A1 (new_n6848_) );
   NAND3_X1 g5393 (
	   .ZN (new_n12124_),
	   .A3 (_net_6958),
	   .A2 (net_6880),
	   .A1 (new_n6846_) );
   NAND2_X1 g5392 (
	   .ZN (new_n12123_),
	   .A2 (net_6848),
	   .A1 (new_n6844_) );
   NAND2_X1 g5391 (
	   .ZN (new_n12122_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n10779_) );
   AND3_X1 g5390 (
	   .ZN (new_n12121_),
	   .A3 (new_n12120_),
	   .A2 (new_n12119_),
	   .A1 (new_n12118_) );
   NAND4_X1 g5389 (
	   .ZN (new_n12120_),
	   .A4 (new_n6841_),
	   .A3 (net_6924),
	   .A2 (_net_6957),
	   .A1 (new_n6829_) );
   NAND4_X1 g5388 (
	   .ZN (new_n12119_),
	   .A4 (new_n6836_1_),
	   .A3 (_net_6957),
	   .A2 (net_6860),
	   .A1 (new_n6838_) );
   NAND4_X1 g5387 (
	   .ZN (new_n12118_),
	   .A4 (new_n6833_),
	   .A3 (_net_6957),
	   .A2 (net_6892),
	   .A1 (new_n6830_) );
   NOR4_X1 g5386 (
	   .ZN (n9709),
	   .A4 (_net_6407),
	   .A3 (new_n9682_),
	   .A2 (new_n9685_),
	   .A1 (new_n10476_) );
   CLKBUF_X1 g5385 (
	   .Z (n9704),
	   .A (_net_7804) );
   NOR2_X1 g5384 (
	   .ZN (n9700),
	   .A2 (new_n12114_),
	   .A1 (new_n12113_) );
   XNOR2_X1 g5383 (
	   .ZN (new_n12114_),
	   .B (new_n12006_),
	   .A (new_n8216_1_) );
   NAND4_X1 g5382 (
	   .ZN (new_n12113_),
	   .A4 (new_n12112_),
	   .A3 (new_n12111_),
	   .A2 (new_n12110_),
	   .A1 (new_n12109_) );
   NAND3_X1 g5381 (
	   .ZN (new_n12112_),
	   .A3 (new_n7135_),
	   .A2 (new_n10008_),
	   .A1 (new_n10418_) );
   NAND2_X1 g5380 (
	   .ZN (new_n12111_),
	   .A2 (_net_6692),
	   .A1 (new_n10419_) );
   NAND2_X1 g5379 (
	   .ZN (new_n12110_),
	   .A2 (new_n6999_),
	   .A1 (new_n7230_1_) );
   OAI21_X1 g5378 (
	   .ZN (new_n12109_),
	   .B2 (new_n6997_),
	   .B1 (n548),
	   .A (_net_6687) );
   CLKBUF_X1 g5377 (
	   .Z (n9695),
	   .A (net_6381) );
   CLKBUF_X1 g5376 (
	   .Z (n9692),
	   .A (net_6703) );
   CLKBUF_X1 g5375 (
	   .Z (n9687),
	   .A (net_6392) );
   MUX2_X1 g5374 (
	   .Z (n9683),
	   .S (new_n10364_),
	   .B (_net_7560),
	   .A (new_n9910_) );
   NOR3_X1 g5373 (
	   .ZN (n9678),
	   .A3 (new_n6891_),
	   .A2 (new_n12103_),
	   .A1 (new_n8958_1_) );
   INV_X1 g5372 (
	   .ZN (new_n12103_),
	   .A (new_n8959_) );
   MUX2_X1 g5371 (
	   .Z (n9673),
	   .S (new_n7028_),
	   .B (_net_7588),
	   .A (new_n8475_) );
   CLKBUF_X1 g5370 (
	   .Z (n9668),
	   .A (net_6383) );
   MUX2_X1 g5369 (
	   .Z (n9664),
	   .S (new_n7544_),
	   .B (_net_7656),
	   .A (new_n9910_) );
   CLKBUF_X1 g5368 (
	   .Z (n9660),
	   .A (net_7005) );
   OAI21_X1 g5367 (
	   .ZN (n9655),
	   .B2 (new_n7222_),
	   .B1 (new_n12097_),
	   .A (new_n12096_) );
   INV_X1 g5366 (
	   .ZN (new_n12097_),
	   .A (_net_7327) );
   NAND2_X1 g5365 (
	   .ZN (new_n12096_),
	   .A2 (new_n8105_),
	   .A1 (new_n7221_1_) );
   CLKBUF_X1 g5364 (
	   .Z (n9651),
	   .A (net_7548) );
   CLKBUF_X1 g5363 (
	   .Z (n9647),
	   .A (net_7386) );
   CLKBUF_X1 g5362 (
	   .Z (n9642),
	   .A (_net_7814) );
   OAI21_X1 g5361 (
	   .ZN (n9638),
	   .B2 (new_n7646_),
	   .B1 (new_n12091_),
	   .A (new_n12090_) );
   INV_X1 g5360 (
	   .ZN (new_n12091_),
	   .A (_net_7414) );
   NAND2_X1 g5359 (
	   .ZN (new_n12090_),
	   .A2 (new_n9037_1_),
	   .A1 (new_n7645_) );
   OAI21_X1 g5358 (
	   .ZN (n9633),
	   .B2 (new_n7272_),
	   .B1 (new_n12088_),
	   .A (new_n12087_) );
   INV_X1 g5357 (
	   .ZN (new_n12088_),
	   .A (_net_7436) );
   NAND2_X1 g5356 (
	   .ZN (new_n12087_),
	   .A2 (new_n8066_),
	   .A1 (new_n7271_) );
   CLKBUF_X1 g5355 (
	   .Z (n9628),
	   .A (net_153) );
   CLKBUF_X1 g5354 (
	   .Z (n9624),
	   .A (_net_7803) );
   CLKBUF_X1 g5353 (
	   .Z (n9620),
	   .A (_net_7820) );
   NOR4_X1 g5352 (
	   .ZN (n9616),
	   .A4 (new_n8186_),
	   .A3 (new_n8185_),
	   .A2 (new_n9685_),
	   .A1 (new_n9844_1_) );
   CLKBUF_X1 g5351 (
	   .Z (n9611),
	   .A (_net_6111) );
   CLKBUF_X1 g5350 (
	   .Z (n9606),
	   .A (_net_7821) );
   OAI21_X1 g5349 (
	   .ZN (n9602),
	   .B2 (new_n7222_),
	   .B1 (new_n12079_),
	   .A (new_n12078_) );
   INV_X1 g5348 (
	   .ZN (new_n12079_),
	   .A (_net_7324) );
   NAND2_X1 g5347 (
	   .ZN (new_n12078_),
	   .A2 (new_n10131_),
	   .A1 (new_n7221_1_) );
   NAND3_X1 g5346 (
	   .ZN (n9597),
	   .A3 (new_n12076_),
	   .A2 (new_n12075_),
	   .A1 (new_n12071_) );
   AOI22_X1 g5345 (
	   .ZN (new_n12076_),
	   .B2 (new_n8180_),
	   .B1 (net_7081),
	   .A2 (new_n7059_),
	   .A1 (new_n10526_) );
   AND3_X1 g5344 (
	   .ZN (new_n12075_),
	   .A3 (new_n12074_),
	   .A2 (new_n12073_),
	   .A1 (new_n12072_) );
   NAND2_X1 g5343 (
	   .ZN (new_n12074_),
	   .A2 (_net_6153),
	   .A1 (new_n7091_) );
   NAND2_X1 g5342 (
	   .ZN (new_n12073_),
	   .A2 (new_n7069_),
	   .A1 (new_n8179_1_) );
   NAND2_X1 g5341 (
	   .ZN (new_n12072_),
	   .A2 (new_n7088_),
	   .A1 (new_n8171_) );
   AND3_X1 g5340 (
	   .ZN (new_n12071_),
	   .A3 (new_n12070_),
	   .A2 (new_n12069_),
	   .A1 (new_n12068_) );
   NAND4_X1 g5339 (
	   .ZN (new_n12070_),
	   .A4 (new_n7044_),
	   .A3 (net_7049),
	   .A2 (_net_7092),
	   .A1 (new_n8154_) );
   NAND4_X1 g5338 (
	   .ZN (new_n12069_),
	   .A4 (new_n7052_),
	   .A3 (net_6985),
	   .A2 (_net_7092),
	   .A1 (new_n8158_) );
   NAND4_X1 g5337 (
	   .ZN (new_n12068_),
	   .A4 (new_n7050_),
	   .A3 (net_7017),
	   .A2 (_net_7092),
	   .A1 (new_n8155_) );
   CLKBUF_X1 g5336 (
	   .Z (n9588),
	   .A (net_6455) );
   OAI21_X1 g5335 (
	   .ZN (n9583),
	   .B2 (new_n7733_),
	   .B1 (new_n9939_1_),
	   .A (new_n12065_) );
   NAND2_X1 g5334 (
	   .ZN (new_n12065_),
	   .A2 (new_n6935_),
	   .A1 (new_n7732_1_) );
   CLKBUF_X1 g5333 (
	   .Z (n9579),
	   .A (net_6840) );
   AOI21_X1 g5332 (
	   .ZN (n9574),
	   .B2 (new_n10248_),
	   .B1 (new_n10247_),
	   .A (new_n8325_) );
   OAI21_X1 g5331 (
	   .ZN (n9569),
	   .B2 (new_n7733_),
	   .B1 (new_n10692_),
	   .A (new_n12061_) );
   NAND2_X1 g5330 (
	   .ZN (new_n12061_),
	   .A2 (new_n8679_),
	   .A1 (new_n7732_1_) );
   MUX2_X1 g5329 (
	   .Z (n9564),
	   .S (new_n7436_),
	   .B (_net_6021),
	   .A (_net_7821) );
   NOR2_X1 g5328 (
	   .ZN (n9559),
	   .A2 (new_n7938_),
	   .A1 (new_n10058_) );
   AOI21_X1 g5327 (
	   .ZN (n9554),
	   .B2 (net_306),
	   .B1 (_net_6018),
	   .A (new_n12057_) );
   NAND3_X1 g5326 (
	   .ZN (new_n12057_),
	   .A3 (_net_6017),
	   .A2 (new_n12056_),
	   .A1 (new_n7655_) );
   INV_X1 g5325 (
	   .ZN (new_n12056_),
	   .A (net_7756) );
   AND2_X1 g5324 (
	   .ZN (n9549),
	   .A2 (net_361),
	   .A1 (new_n6898_) );
   OR4_X1 g5323 (
	   .ZN (n9546),
	   .A4 (new_n12053_),
	   .A3 (new_n12049_),
	   .A2 (new_n12044_),
	   .A1 (new_n12039_) );
   NAND3_X1 g5322 (
	   .ZN (new_n12053_),
	   .A3 (new_n12052_),
	   .A2 (new_n12051_),
	   .A1 (new_n12050_) );
   AOI22_X1 g5321 (
	   .ZN (new_n12052_),
	   .B2 (_net_7700),
	   .B1 (_net_7729),
	   .A2 (_net_7723),
	   .A1 (_net_7694) );
   AOI22_X1 g5320 (
	   .ZN (new_n12051_),
	   .B2 (_net_7695),
	   .B1 (_net_7724),
	   .A2 (_net_7701),
	   .A1 (_net_7730) );
   AOI22_X1 g5319 (
	   .ZN (new_n12050_),
	   .B2 (_net_7745),
	   .B1 (_net_7716),
	   .A2 (_net_7705),
	   .A1 (_net_7734) );
   NAND4_X1 g5318 (
	   .ZN (new_n12049_),
	   .A4 (new_n12048_),
	   .A3 (new_n12047_),
	   .A2 (new_n12046_),
	   .A1 (new_n12045_) );
   NAND2_X1 g5317 (
	   .ZN (new_n12048_),
	   .A2 (_net_7733),
	   .A1 (_net_7704) );
   AOI22_X1 g5316 (
	   .ZN (new_n12047_),
	   .B2 (net_7712),
	   .B1 (net_7741),
	   .A2 (net_7709),
	   .A1 (net_7738) );
   AOI22_X1 g5315 (
	   .ZN (new_n12046_),
	   .B2 (net_7739),
	   .B1 (net_7710),
	   .A2 (net_7737),
	   .A1 (net_7708) );
   AOI22_X1 g5314 (
	   .ZN (new_n12045_),
	   .B2 (net_7715),
	   .B1 (net_7744),
	   .A2 (net_7714),
	   .A1 (net_7743) );
   NAND4_X1 g5313 (
	   .ZN (new_n12044_),
	   .A4 (new_n12043_),
	   .A3 (new_n12042_),
	   .A2 (new_n12041_),
	   .A1 (new_n12040_) );
   AOI22_X1 g5312 (
	   .ZN (new_n12043_),
	   .B2 (_net_7721),
	   .B1 (_net_7692),
	   .A2 (_net_7719),
	   .A1 (_net_7748) );
   AOI22_X1 g5311 (
	   .ZN (new_n12042_),
	   .B2 (_net_7699),
	   .B1 (_net_7728),
	   .A2 (_net_7725),
	   .A1 (_net_7696) );
   AOI22_X1 g5310 (
	   .ZN (new_n12041_),
	   .B2 (_net_7726),
	   .B1 (_net_7697),
	   .A2 (_net_7736),
	   .A1 (_net_7707) );
   AOI22_X1 g5309 (
	   .ZN (new_n12040_),
	   .B2 (_net_7693),
	   .B1 (_net_7722),
	   .A2 (net_7742),
	   .A1 (net_7713) );
   NAND4_X1 g5308 (
	   .ZN (new_n12039_),
	   .A4 (new_n12038_),
	   .A3 (new_n12037_),
	   .A2 (new_n12036_),
	   .A1 (new_n12035_) );
   AOI22_X1 g5307 (
	   .ZN (new_n12038_),
	   .B2 (_net_7735),
	   .B1 (_net_7706),
	   .A2 (net_7691),
	   .A1 (_net_7720) );
   AOI22_X1 g5306 (
	   .ZN (new_n12037_),
	   .B2 (_net_7702),
	   .B1 (_net_7731),
	   .A2 (_net_7703),
	   .A1 (_net_7732) );
   AOI22_X1 g5305 (
	   .ZN (new_n12036_),
	   .B2 (net_7740),
	   .B1 (net_7711),
	   .A2 (_net_7718),
	   .A1 (_net_7747) );
   AOI22_X1 g5304 (
	   .ZN (new_n12035_),
	   .B2 (_net_7727),
	   .B1 (_net_7698),
	   .A2 (_net_7717),
	   .A1 (_net_7746) );
   CLKBUF_X1 g5303 (
	   .Z (n9541),
	   .A (_net_7813) );
   CLKBUF_X1 g5302 (
	   .Z (n9537),
	   .A (_net_7817) );
   NAND2_X1 g5301 (
	   .ZN (n9533),
	   .A2 (new_n12031_),
	   .A1 (new_n12030_) );
   AOI22_X1 g5300 (
	   .ZN (new_n12031_),
	   .B2 (net_7521),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7489) );
   AOI22_X1 g5299 (
	   .ZN (new_n12030_),
	   .B2 (_net_7425),
	   .B1 (new_n7298_),
	   .A2 (net_7457),
	   .A1 (new_n7296_) );
   CLKBUF_X1 g5298 (
	   .Z (n9528),
	   .A (_net_7805) );
   CLKBUF_X1 g5297 (
	   .Z (n9525),
	   .A (net_7015) );
   CLKBUF_X1 g5296 (
	   .Z (n9520),
	   .A (net_6391) );
   CLKBUF_X1 g5295 (
	   .Z (n9517),
	   .A (net_6871) );
   MUX2_X1 g5294 (
	   .Z (n9512),
	   .S (new_n7503_),
	   .B (_net_7616),
	   .A (new_n8899_1_) );
   MUX2_X1 g5293 (
	   .Z (n9507),
	   .S (new_n7503_),
	   .B (_net_7617),
	   .A (new_n8336_) );
   CLKBUF_X1 g5292 (
	   .Z (n9502),
	   .A (_net_6163) );
   MUX2_X1 g5291 (
	   .Z (n9497),
	   .S (new_n7028_),
	   .B (_net_7597),
	   .A (new_n7523_) );
   OAI21_X1 g5290 (
	   .ZN (n9492),
	   .B2 (new_n7252_1_),
	   .B1 (new_n10673_),
	   .A (new_n12020_) );
   NAND2_X1 g5289 (
	   .ZN (new_n12020_),
	   .A2 (new_n8780_1_),
	   .A1 (new_n7251_) );
   OAI21_X1 g5288 (
	   .ZN (n9487),
	   .B2 (new_n7646_),
	   .B1 (new_n12018_),
	   .A (new_n12017_) );
   INV_X1 g5287 (
	   .ZN (new_n12018_),
	   .A (_net_7415) );
   NAND2_X1 g5286 (
	   .ZN (new_n12017_),
	   .A2 (new_n7595_),
	   .A1 (new_n7645_) );
   CLKBUF_X1 g5285 (
	   .Z (n9483),
	   .A (net_6611) );
   NOR2_X1 g5284 (
	   .ZN (n9478),
	   .A2 (new_n9900_),
	   .A1 (new_n7035_) );
   CLKBUF_X1 g5283 (
	   .Z (n9475),
	   .A (net_6842) );
   CLKBUF_X1 g5282 (
	   .Z (n9470),
	   .A (net_6394) );
   CLKBUF_X1 g5281 (
	   .Z (n9467),
	   .A (net_6972) );
   CLKBUF_X1 g5280 (
	   .Z (n9462),
	   .A (_net_7816) );
   CLKBUF_X1 g5279 (
	   .Z (n9459),
	   .A (net_7709) );
   OAI21_X1 g5278 (
	   .ZN (n9454),
	   .B2 (new_n12008_),
	   .B1 (new_n12004_),
	   .A (new_n10006_1_) );
   OAI21_X1 g5277 (
	   .ZN (new_n12008_),
	   .B2 (new_n12007_),
	   .B1 (new_n12005_),
	   .A (new_n7779_1_) );
   NOR2_X1 g5276 (
	   .ZN (new_n12007_),
	   .A2 (_net_6690),
	   .A1 (new_n12006_) );
   INV_X1 g5275 (
	   .ZN (new_n12006_),
	   .A (_net_6693) );
   NOR2_X1 g5274 (
	   .ZN (new_n12005_),
	   .A2 (_net_6693),
	   .A1 (new_n8214_) );
   NAND2_X1 g5273 (
	   .ZN (new_n12004_),
	   .A2 (_net_5967),
	   .A1 (n548) );
   AND2_X1 g5272 (
	   .ZN (n9449),
	   .A2 (_net_6319),
	   .A1 (new_n7235_1_) );
   CLKBUF_X1 g5271 (
	   .Z (n9445),
	   .A (net_6731) );
   NAND4_X1 g5270 (
	   .ZN (n9441),
	   .A4 (new_n12000_),
	   .A3 (new_n11999_),
	   .A2 (new_n11998_),
	   .A1 (new_n11997_) );
   NAND4_X1 g5269 (
	   .ZN (new_n12000_),
	   .A4 (new_n7364_),
	   .A3 (_net_5991),
	   .A2 (x1322),
	   .A1 (new_n7399_) );
   NAND4_X1 g5268 (
	   .ZN (new_n11999_),
	   .A4 (_net_7698),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   NAND4_X1 g5267 (
	   .ZN (new_n11998_),
	   .A4 (net_274),
	   .A3 (x1286),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR2_X1 g5266 (
	   .ZN (new_n11997_),
	   .A2 (new_n11996_),
	   .A1 (new_n11991_) );
   NAND4_X1 g5265 (
	   .ZN (new_n11996_),
	   .A4 (new_n11995_),
	   .A3 (new_n11994_),
	   .A2 (new_n11993_),
	   .A1 (new_n11992_) );
   NAND4_X1 g5264 (
	   .ZN (new_n11995_),
	   .A4 (net_163),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g5263 (
	   .ZN (new_n11994_),
	   .A3 (net_200),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g5262 (
	   .ZN (new_n11993_),
	   .A3 (net_237),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   NAND4_X1 g5261 (
	   .ZN (new_n11992_),
	   .A4 (_net_7727),
	   .A3 (x1286),
	   .A2 (x1261),
	   .A1 (new_n7370_) );
   NAND2_X1 g5260 (
	   .ZN (new_n11991_),
	   .A2 (new_n11990_),
	   .A1 (new_n11989_) );
   NAND4_X1 g5259 (
	   .ZN (new_n11990_),
	   .A4 (new_n7354_1_),
	   .A3 (_net_121),
	   .A2 (x1261),
	   .A1 (new_n7370_) );
   NAND4_X1 g5258 (
	   .ZN (new_n11989_),
	   .A4 (new_n7371_),
	   .A3 (new_n7370_),
	   .A2 (net_6035),
	   .A1 (new_n7369_) );
   AOI21_X1 g5257 (
	   .ZN (n9436),
	   .B2 (new_n11987_),
	   .B1 (new_n11842_),
	   .A (new_n7427_1_) );
   INV_X1 g5256 (
	   .ZN (new_n11987_),
	   .A (_net_288) );
   CLKBUF_X1 g5255 (
	   .Z (n9431),
	   .A (_net_7810) );
   CLKBUF_X1 g5254 (
	   .Z (n9428),
	   .A (_net_7808) );
   CLKBUF_X1 g5253 (
	   .Z (n9425),
	   .A (net_6459) );
   OAI21_X1 g5252 (
	   .ZN (n9420),
	   .B2 (new_n7222_),
	   .B1 (new_n11982_),
	   .A (new_n11981_) );
   INV_X1 g5251 (
	   .ZN (new_n11982_),
	   .A (_net_7317) );
   NAND2_X1 g5250 (
	   .ZN (new_n11981_),
	   .A2 (new_n7255_),
	   .A1 (new_n7221_1_) );
   OAI21_X1 g5249 (
	   .ZN (n9415),
	   .B2 (new_n10086_),
	   .B1 (new_n11979_),
	   .A (new_n11978_) );
   INV_X1 g5248 (
	   .ZN (new_n11979_),
	   .A (_net_6085) );
   NAND2_X1 g5247 (
	   .ZN (new_n11978_),
	   .A2 (new_n6980_),
	   .A1 (new_n8123_) );
   MUX2_X1 g5246 (
	   .Z (n9410),
	   .S (new_n10364_),
	   .B (_net_7569),
	   .A (new_n9349_) );
   CLKBUF_X1 g5245 (
	   .Z (n9405),
	   .A (_net_7808) );
   CLKBUF_X1 g5244 (
	   .Z (n9402),
	   .A (x0) );
   CLKBUF_X1 g5243 (
	   .Z (n9398),
	   .A (_net_6102) );
   CLKBUF_X1 g5242 (
	   .Z (n9393),
	   .A (_net_7804) );
   CLKBUF_X1 g5241 (
	   .Z (n9390),
	   .A (net_6601) );
   CLKBUF_X1 g5240 (
	   .Z (n9385),
	   .A (_net_7805) );
   CLKBUF_X1 g5239 (
	   .Z (n9381),
	   .A (_net_7821) );
   CLKBUF_X1 g5238 (
	   .Z (n9377),
	   .A (_net_7820) );
   CLKBUF_X1 g5237 (
	   .Z (n9373),
	   .A (_net_7810) );
   CLKBUF_X1 g5236 (
	   .Z (n9370),
	   .A (net_7099) );
   CLKBUF_X1 g5235 (
	   .Z (n9365),
	   .A (_net_6089) );
   CLKBUF_X1 g5234 (
	   .Z (n9361),
	   .A (net_6464) );
   CLKBUF_X1 g5233 (
	   .Z (n9356),
	   .A (_net_7794) );
   OAI21_X1 g5232 (
	   .ZN (n9352),
	   .B2 (new_n7733_),
	   .B1 (new_n11364_),
	   .A (new_n11962_) );
   NAND2_X1 g5231 (
	   .ZN (new_n11962_),
	   .A2 (new_n8229_),
	   .A1 (new_n7732_1_) );
   CLKBUF_X1 g5230 (
	   .Z (n9348),
	   .A (net_7541) );
   CLKBUF_X1 g5229 (
	   .Z (n9343),
	   .A (_net_7808) );
   CLKBUF_X1 g5228 (
	   .Z (n9339),
	   .A (_net_7800) );
   AOI21_X1 g5227 (
	   .ZN (n9335),
	   .B2 (new_n10798_),
	   .B1 (new_n11957_),
	   .A (new_n7427_1_) );
   INV_X1 g5226 (
	   .ZN (new_n11957_),
	   .A (net_6003) );
   NOR2_X1 g5225 (
	   .ZN (n9330),
	   .A2 (new_n7878_1_),
	   .A1 (new_n9927_) );
   CLKBUF_X1 g5224 (
	   .Z (n9326),
	   .A (net_6749) );
   NAND2_X1 g5223 (
	   .ZN (n9321),
	   .A2 (new_n11953_),
	   .A1 (new_n11952_) );
   AOI22_X1 g5222 (
	   .ZN (new_n11953_),
	   .B2 (net_7523),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7491) );
   AOI22_X1 g5221 (
	   .ZN (new_n11952_),
	   .B2 (_net_7427),
	   .B1 (new_n7298_),
	   .A2 (net_7459),
	   .A1 (new_n7296_) );
   NOR2_X1 g5220 (
	   .ZN (n9316),
	   .A2 (new_n7602_),
	   .A1 (new_n8675_) );
   AOI21_X1 g5219 (
	   .ZN (n9312),
	   .B2 (new_n7619_),
	   .B1 (new_n7265_1_),
	   .A (new_n7427_1_) );
   OAI21_X1 g5218 (
	   .ZN (n9307),
	   .B2 (new_n7733_),
	   .B1 (new_n7304_),
	   .A (new_n11948_) );
   NAND2_X1 g5217 (
	   .ZN (new_n11948_),
	   .A2 (new_n9901_),
	   .A1 (new_n7732_1_) );
   NOR2_X1 g5216 (
	   .ZN (n9302),
	   .A2 (new_n7274_),
	   .A1 (new_n7035_) );
   AND2_X1 g5215 (
	   .ZN (n9298),
	   .A2 (net_382),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g5214 (
	   .Z (n9294),
	   .A (_net_7816) );
   CLKBUF_X1 g5213 (
	   .Z (n9290),
	   .A (_net_7820) );
   CLKBUF_X1 g5212 (
	   .Z (n9287),
	   .A (net_6848) );
   NAND3_X1 g5211 (
	   .ZN (n9282),
	   .A3 (new_n11941_),
	   .A2 (new_n11940_),
	   .A1 (new_n11936_) );
   AOI22_X1 g5210 (
	   .ZN (new_n11941_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6950),
	   .A2 (new_n6851_),
	   .A1 (new_n6879_) );
   AND3_X1 g5209 (
	   .ZN (new_n11940_),
	   .A3 (new_n11939_),
	   .A2 (new_n11938_),
	   .A1 (new_n11937_) );
   NAND2_X1 g5208 (
	   .ZN (new_n11939_),
	   .A2 (_net_6137),
	   .A1 (new_n6868_) );
   NAND2_X1 g5207 (
	   .ZN (new_n11938_),
	   .A2 (new_n6862_),
	   .A1 (new_n7716_) );
   NAND2_X1 g5206 (
	   .ZN (new_n11937_),
	   .A2 (new_n6853_),
	   .A1 (new_n8457_) );
   AND3_X1 g5205 (
	   .ZN (new_n11936_),
	   .A3 (new_n11935_),
	   .A2 (new_n11934_),
	   .A1 (new_n11933_) );
   NAND4_X1 g5204 (
	   .ZN (new_n11935_),
	   .A4 (new_n6841_),
	   .A3 (_net_6957),
	   .A2 (net_6918),
	   .A1 (new_n6829_) );
   NAND4_X1 g5203 (
	   .ZN (new_n11934_),
	   .A4 (new_n6836_1_),
	   .A3 (_net_6957),
	   .A2 (net_6854),
	   .A1 (new_n6838_) );
   NAND4_X1 g5202 (
	   .ZN (new_n11933_),
	   .A4 (new_n6833_),
	   .A3 (_net_6957),
	   .A2 (net_6886),
	   .A1 (new_n6830_) );
   NAND2_X1 g5201 (
	   .ZN (n9277),
	   .A2 (new_n11931_),
	   .A1 (new_n11930_) );
   NAND2_X1 g5200 (
	   .ZN (new_n11931_),
	   .A2 (new_n7587_),
	   .A1 (new_n7198_) );
   AOI22_X1 g5199 (
	   .ZN (new_n11930_),
	   .B2 (new_n7210_),
	   .B1 (_net_6106),
	   .A2 (new_n7203_1_),
	   .A1 (new_n8245_1_) );
   NAND2_X1 g5198 (
	   .ZN (n9272),
	   .A2 (new_n11928_),
	   .A1 (new_n11927_) );
   NAND3_X1 g5197 (
	   .ZN (new_n11928_),
	   .A3 (_net_7530),
	   .A2 (_net_278),
	   .A1 (new_n10359_) );
   OAI21_X1 g5196 (
	   .ZN (new_n11927_),
	   .B2 (new_n7301_),
	   .B1 (new_n7296_),
	   .A (n5792) );
   CLKBUF_X1 g5195 (
	   .Z (n9267),
	   .A (net_7807) );
   OAI21_X1 g5194 (
	   .ZN (n9263),
	   .B2 (new_n7736_),
	   .B1 (new_n9211_1_),
	   .A (new_n11924_) );
   NAND2_X1 g5193 (
	   .ZN (new_n11924_),
	   .A2 (new_n8280_1_),
	   .A1 (new_n7732_1_) );
   OAI21_X1 g5192 (
	   .ZN (n9258),
	   .B2 (new_n11922_),
	   .B1 (new_n9933_),
	   .A (new_n6963_) );
   NOR2_X1 g5191 (
	   .ZN (new_n11922_),
	   .A2 (_net_6405),
	   .A1 (_net_6404) );
   CLKBUF_X1 g5190 (
	   .Z (n9254),
	   .A (net_7103) );
   CLKBUF_X1 g5189 (
	   .Z (n9250),
	   .A (net_6701) );
   CLKBUF_X1 g5188 (
	   .Z (n9245),
	   .A (_net_7800) );
   CLKBUF_X1 g5187 (
	   .Z (n9242),
	   .A (net_6483) );
   CLKBUF_X1 g5186 (
	   .Z (n9238),
	   .A (net_6705) );
   MUX2_X1 g5185 (
	   .Z (n9233),
	   .S (new_n7284_1_),
	   .B (_net_7701),
	   .A (_net_7803) );
   NOR2_X1 g5184 (
	   .ZN (n9228),
	   .A2 (new_n6903_),
	   .A1 (new_n7035_) );
   CLKBUF_X1 g5183 (
	   .Z (n9225),
	   .A (net_7156) );
   NAND3_X1 g5182 (
	   .ZN (n9220),
	   .A3 (new_n11912_),
	   .A2 (new_n11911_),
	   .A1 (new_n11907_) );
   AOI22_X1 g5181 (
	   .ZN (new_n11912_),
	   .B2 (new_n7136_),
	   .B1 (net_6677),
	   .A2 (new_n8939_1_),
	   .A1 (new_n7013_1_) );
   AND3_X1 g5180 (
	   .ZN (new_n11911_),
	   .A3 (new_n11910_),
	   .A2 (new_n11909_),
	   .A1 (new_n11908_) );
   NAND2_X1 g5179 (
	   .ZN (new_n11910_),
	   .A2 (_net_6094),
	   .A1 (new_n6984_) );
   NAND2_X1 g5178 (
	   .ZN (new_n11909_),
	   .A2 (new_n6994_),
	   .A1 (new_n9328_) );
   NAND2_X1 g5177 (
	   .ZN (new_n11908_),
	   .A2 (new_n6979_),
	   .A1 (new_n10181_) );
   AND3_X1 g5176 (
	   .ZN (new_n11907_),
	   .A3 (new_n11906_),
	   .A2 (new_n11905_),
	   .A1 (new_n11904_) );
   NAND4_X1 g5175 (
	   .ZN (new_n11906_),
	   .A4 (new_n6987_),
	   .A3 (net_6645),
	   .A2 (_net_6687),
	   .A1 (new_n7114_) );
   NAND4_X1 g5174 (
	   .ZN (new_n11905_),
	   .A4 (new_n6990_1_),
	   .A3 (net_6581),
	   .A2 (_net_6687),
	   .A1 (new_n7118_) );
   NAND4_X1 g5173 (
	   .ZN (new_n11904_),
	   .A4 (new_n6989_),
	   .A3 (net_6613),
	   .A2 (_net_6687),
	   .A1 (new_n7115_) );
   NOR2_X1 g5172 (
	   .ZN (n9215),
	   .A2 (new_n7107_1_),
	   .A1 (new_n8675_) );
   NOR2_X1 g5171 (
	   .ZN (n9211),
	   .A2 (x940),
	   .A1 (new_n11901_) );
   NAND2_X1 g5170 (
	   .ZN (new_n11901_),
	   .A2 (_net_6034),
	   .A1 (n9592) );
   MUX2_X1 g5169 (
	   .Z (n9206),
	   .S (new_n7436_),
	   .B (_net_5986),
	   .A (_net_7795) );
   AOI21_X1 g5168 (
	   .ZN (n9201),
	   .B2 (new_n10505_),
	   .B1 (_net_7682),
	   .A (new_n11898_) );
   OAI21_X1 g5167 (
	   .ZN (new_n11898_),
	   .B2 (_net_7682),
	   .B1 (new_n10505_),
	   .A (_net_289) );
   CLKBUF_X1 g5166 (
	   .Z (n9196),
	   .A (net_6383) );
   OAI221_X1 g5165 (
	   .ZN (n9192),
	   .C2 (new_n6917_),
	   .C1 (new_n10986_),
	   .B2 (new_n7986_),
	   .B1 (new_n9262_),
	   .A (new_n11895_) );
   AOI22_X1 g5164 (
	   .ZN (new_n11895_),
	   .B2 (_net_7266),
	   .B1 (new_n10556_),
	   .A2 (_net_7330),
	   .A1 (new_n10555_) );
   OAI21_X1 g5163 (
	   .ZN (n9187),
	   .B2 (new_n6949_),
	   .B1 (new_n11893_),
	   .A (new_n11892_) );
   INV_X1 g5162 (
	   .ZN (new_n11893_),
	   .A (_net_7260) );
   NAND2_X1 g5161 (
	   .ZN (new_n11892_),
	   .A2 (new_n10131_),
	   .A1 (new_n6948_) );
   CLKBUF_X1 g5160 (
	   .Z (n9182),
	   .A (_net_7797) );
   CLKBUF_X1 g5159 (
	   .Z (n9178),
	   .A (_net_6077) );
   AND2_X1 g5158 (
	   .ZN (n9173),
	   .A2 (_net_6187),
	   .A1 (new_n7235_1_) );
   CLKBUF_X1 g5157 (
	   .Z (n9169),
	   .A (net_6565) );
   CLKBUF_X1 g5156 (
	   .Z (n9164),
	   .A (_net_7811) );
   CLKBUF_X1 g5155 (
	   .Z (n9160),
	   .A (net_6393) );
   OAI21_X1 g5154 (
	   .ZN (n9156),
	   .B2 (new_n6949_),
	   .B1 (new_n11884_),
	   .A (new_n11883_) );
   INV_X1 g5153 (
	   .ZN (new_n11884_),
	   .A (_net_7259) );
   NAND2_X1 g5152 (
	   .ZN (new_n11883_),
	   .A2 (new_n7108_),
	   .A1 (new_n6948_) );
   OAI221_X1 g5151 (
	   .ZN (n9151),
	   .C2 (new_n7312_1_),
	   .C1 (new_n9839_),
	   .B2 (new_n7986_),
	   .B1 (new_n8294_1_),
	   .A (new_n11881_) );
   AOI22_X1 g5150 (
	   .ZN (new_n11881_),
	   .B2 (_net_7256),
	   .B1 (new_n10556_),
	   .A2 (_net_7320),
	   .A1 (new_n10555_) );
   CLKBUF_X1 g5149 (
	   .Z (n9146),
	   .A (_net_7803) );
   CLKBUF_X1 g5148 (
	   .Z (n9143),
	   .A (net_6876) );
   CLKBUF_X1 g5147 (
	   .Z (n9138),
	   .A (_net_7793) );
   CLKBUF_X1 g5146 (
	   .Z (n9134),
	   .A (_net_6137) );
   MUX2_X1 g5145 (
	   .Z (n9129),
	   .S (new_n7544_),
	   .B (_net_7660),
	   .A (new_n8151_) );
   MUX2_X1 g5144 (
	   .Z (n9124),
	   .S (new_n10364_),
	   .B (_net_7558),
	   .A (new_n7762_) );
   CLKBUF_X1 g5143 (
	   .Z (n9120),
	   .A (net_7155) );
   MUX2_X1 g5142 (
	   .Z (n9115),
	   .S (new_n7537_),
	   .B (_net_292),
	   .A (_net_7812) );
   CLKBUF_X1 g5141 (
	   .Z (n9110),
	   .A (x1511) );
   MUX2_X1 g5140 (
	   .Z (n9106),
	   .S (new_n7284_1_),
	   .B (_net_7716),
	   .A (_net_7818) );
   MUX2_X1 g5139 (
	   .Z (n9101),
	   .S (new_n7537_),
	   .B (_net_289),
	   .A (_net_7809) );
   NAND2_X1 g5138 (
	   .ZN (n9096),
	   .A2 (new_n11868_),
	   .A1 (new_n11867_) );
   AOI22_X1 g5137 (
	   .ZN (new_n11868_),
	   .B2 (_net_7578),
	   .B1 (new_n6751_),
	   .A2 (net_7610),
	   .A1 (new_n6743_) );
   AOI22_X1 g5136 (
	   .ZN (new_n11867_),
	   .B2 (net_7642),
	   .B1 (new_n8009_),
	   .A2 (new_n7970_1_),
	   .A1 (net_7674) );
   CLKBUF_X1 g5135 (
	   .Z (n9091),
	   .A (_net_6094) );
   CLKBUF_X1 g5134 (
	   .Z (n9086),
	   .A (_net_7819) );
   CLKBUF_X1 g5133 (
	   .Z (n9082),
	   .A (_net_7817) );
   CLKBUF_X1 g5132 (
	   .Z (n9079),
	   .A (net_7101) );
   MUX2_X1 g5131 (
	   .Z (n9074),
	   .S (_net_154),
	   .B (net_311),
	   .A (_net_115) );
   CLKBUF_X1 g5130 (
	   .Z (n9069),
	   .A (_net_6110) );
   CLKBUF_X1 g5129 (
	   .Z (n9065),
	   .A (net_6984) );
   NOR2_X1 g5128 (
	   .ZN (n9060),
	   .A2 (new_n7104_),
	   .A1 (new_n8675_) );
   CLKBUF_X1 g5127 (
	   .Z (n9057),
	   .A (net_6966) );
   AOI21_X1 g5126 (
	   .ZN (n9052),
	   .B2 (new_n7739_),
	   .B1 (new_n11856_),
	   .A (new_n11855_) );
   INV_X1 g5125 (
	   .ZN (new_n11856_),
	   .A (_net_7423) );
   NOR2_X1 g5124 (
	   .ZN (new_n11855_),
	   .A2 (n634),
	   .A1 (new_n7738_) );
   CLKBUF_X1 g5123 (
	   .Z (n9047),
	   .A (_net_189) );
   NAND2_X1 g5122 (
	   .ZN (n9042),
	   .A2 (new_n11852_),
	   .A1 (new_n11851_) );
   AOI22_X1 g5121 (
	   .ZN (new_n11852_),
	   .B2 (_net_7552),
	   .B1 (new_n6751_),
	   .A2 (_net_7616),
	   .A1 (new_n6746_1_) );
   AOI22_X1 g5120 (
	   .ZN (new_n11851_),
	   .B2 (_net_7584),
	   .B1 (new_n7350_),
	   .A2 (new_n7970_1_),
	   .A1 (_net_7648) );
   CLKBUF_X1 g5119 (
	   .Z (n9037),
	   .A (_net_7805) );
   CLKBUF_X1 g5118 (
	   .Z (n9034),
	   .A (net_6864) );
   OAI211_X1 g5117 (
	   .ZN (n9030),
	   .C2 (new_n7366_),
	   .C1 (new_n11847_),
	   .B (new_n11846_),
	   .A (new_n11845_) );
   INV_X1 g5116 (
	   .ZN (new_n11847_),
	   .A (_net_6018) );
   NAND4_X1 g5115 (
	   .ZN (new_n11846_),
	   .A4 (_net_7716),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   NOR3_X1 g5114 (
	   .ZN (new_n11845_),
	   .A3 (new_n11844_),
	   .A2 (new_n11843_),
	   .A1 (new_n11841_) );
   AND3_X1 g5113 (
	   .ZN (new_n11844_),
	   .A3 (new_n7382_),
	   .A2 (net_255),
	   .A1 (new_n7380_) );
   NOR2_X1 g5112 (
	   .ZN (new_n11843_),
	   .A2 (new_n11842_),
	   .A1 (new_n7378_) );
   INV_X1 g5111 (
	   .ZN (new_n11842_),
	   .A (_net_7745) );
   OAI22_X1 g5110 (
	   .ZN (new_n11841_),
	   .B2 (new_n11840_),
	   .B1 (new_n7938_),
	   .A2 (new_n11839_),
	   .A1 (new_n7936_) );
   INV_X1 g5109 (
	   .ZN (new_n11840_),
	   .A (net_181) );
   INV_X1 g5108 (
	   .ZN (new_n11839_),
	   .A (net_218) );
   CLKBUF_X1 g5107 (
	   .Z (n9025),
	   .A (_net_7800) );
   CLKBUF_X1 g5106 (
	   .Z (n9022),
	   .A (net_6445) );
   CLKBUF_X1 g5105 (
	   .Z (n9017),
	   .A (net_136) );
   CLKBUF_X1 g5104 (
	   .Z (n9014),
	   .A (net_7017) );
   CLKBUF_X1 g5103 (
	   .Z (n9010),
	   .A (net_6582) );
   OAI21_X1 g5102 (
	   .ZN (n9005),
	   .B2 (new_n11832_),
	   .B1 (new_n9345_),
	   .A (new_n11831_) );
   OR2_X1 g5101 (
	   .ZN (new_n11832_),
	   .A2 (_net_7783),
	   .A1 (new_n9950_) );
   OAI211_X1 g5100 (
	   .ZN (new_n11831_),
	   .C2 (new_n9950_),
	   .C1 (new_n9341_),
	   .B (_net_7783),
	   .A (new_n9342_) );
   OAI21_X1 g5099 (
	   .ZN (n9000),
	   .B2 (new_n7538_),
	   .B1 (new_n8091_),
	   .A (new_n11829_) );
   NAND2_X1 g5098 (
	   .ZN (new_n11829_),
	   .A2 (_net_268),
	   .A1 (new_n7538_) );
   MUX2_X1 g5097 (
	   .Z (n8995),
	   .S (new_n7537_),
	   .B (_net_293),
	   .A (_net_7813) );
   CLKBUF_X1 g5096 (
	   .Z (n8990),
	   .A (net_6386) );
   MUX2_X1 g5095 (
	   .Z (n8986),
	   .S (new_n10364_),
	   .B (_net_7581),
	   .A (n698) );
   CLKBUF_X1 g5094 (
	   .Z (n8981),
	   .A (_net_6154) );
   OAI21_X1 g5093 (
	   .ZN (n8976),
	   .B2 (new_n6897_),
	   .B1 (new_n10955_),
	   .A (new_n11823_) );
   NAND2_X1 g5092 (
	   .ZN (new_n11823_),
	   .A2 (new_n7991_),
	   .A1 (new_n6896_) );
   CLKBUF_X1 g5091 (
	   .Z (n8971),
	   .A (net_7807) );
   OAI221_X1 g5090 (
	   .ZN (n8967),
	   .C2 (new_n7306_),
	   .C1 (new_n10216_),
	   .B2 (new_n7302_1_),
	   .B1 (new_n6906_1_),
	   .A (new_n11820_) );
   AOI22_X1 g5089 (
	   .ZN (new_n11820_),
	   .B2 (_net_7417),
	   .B1 (new_n9203_),
	   .A2 (_net_7449),
	   .A1 (new_n7295_) );
   CLKBUF_X1 g5088 (
	   .Z (n8963),
	   .A (net_7544) );
   CLKBUF_X1 g5087 (
	   .Z (n8958),
	   .A (_net_6130) );
   OAI21_X1 g5086 (
	   .ZN (n8953),
	   .B2 (new_n7272_),
	   .B1 (new_n11816_),
	   .A (new_n11815_) );
   INV_X1 g5085 (
	   .ZN (new_n11816_),
	   .A (_net_7451) );
   NAND2_X1 g5084 (
	   .ZN (new_n11815_),
	   .A2 (new_n8280_1_),
	   .A1 (new_n7271_) );
   OAI21_X1 g5083 (
	   .ZN (n8948),
	   .B2 (new_n7222_),
	   .B1 (new_n11813_),
	   .A (new_n11812_) );
   INV_X1 g5082 (
	   .ZN (new_n11813_),
	   .A (_net_7322) );
   NAND2_X1 g5081 (
	   .ZN (new_n11812_),
	   .A2 (new_n7495_),
	   .A1 (new_n7221_1_) );
   CLKBUF_X1 g5080 (
	   .Z (n8943),
	   .A (_net_6086) );
   CLKBUF_X1 g5079 (
	   .Z (n8939),
	   .A (net_6458) );
   NOR2_X1 g5078 (
	   .ZN (n8934),
	   .A2 (new_n7494_),
	   .A1 (new_n8675_) );
   CLKBUF_X1 g5077 (
	   .Z (n8931),
	   .A (net_7243) );
   CLKBUF_X1 g5076 (
	   .Z (n8926),
	   .A (_net_7809) );
   NOR3_X1 g5075 (
	   .ZN (n8922),
	   .A3 (new_n11805_),
	   .A2 (new_n10597_),
	   .A1 (new_n7449_) );
   NOR2_X1 g5074 (
	   .ZN (new_n11805_),
	   .A2 (_net_7787),
	   .A1 (new_n7451_) );
   NAND2_X1 g5073 (
	   .ZN (n8917),
	   .A2 (new_n11803_),
	   .A1 (new_n11802_) );
   NAND2_X1 g5072 (
	   .ZN (new_n11803_),
	   .A2 (new_n7701_),
	   .A1 (new_n8034_) );
   AOI22_X1 g5071 (
	   .ZN (new_n11802_),
	   .B2 (new_n7694_),
	   .B1 (_net_6166),
	   .A2 (new_n7690_),
	   .A1 (new_n8030_) );
   CLKBUF_X1 g5070 (
	   .Z (n8912),
	   .A (_net_7804) );
   CLKBUF_X1 g5069 (
	   .Z (n8908),
	   .A (_net_6119) );
   CLKBUF_X1 g5068 (
	   .Z (n8903),
	   .A (_net_7822) );
   NOR2_X1 g5067 (
	   .ZN (n8899),
	   .A2 (new_n7493_),
	   .A1 (new_n8675_) );
   AND2_X1 g5066 (
	   .ZN (n8895),
	   .A2 (_net_6297),
	   .A1 (new_n7235_1_) );
   CLKBUF_X1 g5065 (
	   .Z (n8891),
	   .A (net_7132) );
   CLKBUF_X1 g5064 (
	   .Z (n8886),
	   .A (_net_7819) );
   CLKBUF_X1 g5063 (
	   .Z (n8882),
	   .A (net_6060) );
   CLKBUF_X1 g5062 (
	   .Z (n8877),
	   .A (net_6389) );
   CLKBUF_X1 g5061 (
	   .Z (n8873),
	   .A (net_151) );
   AND2_X1 g5060 (
	   .ZN (n8869),
	   .A2 (_net_6185),
	   .A1 (new_n7235_1_) );
   CLKBUF_X1 g5059 (
	   .Z (n8864),
	   .A (x1494) );
   MUX2_X1 g5058 (
	   .Z (n8860),
	   .S (new_n7503_),
	   .B (_net_7625),
	   .A (new_n10112_1_) );
   OAI21_X1 g5057 (
	   .ZN (n8855),
	   .B2 (new_n7101_),
	   .B1 (new_n8948_1_),
	   .A (new_n11787_) );
   NAND2_X1 g5056 (
	   .ZN (new_n11787_),
	   .A2 (new_n7667_),
	   .A1 (new_n7100_) );
   OAI21_X1 g5055 (
	   .ZN (n8845),
	   .B2 (new_n11785_),
	   .B1 (new_n7691_1_),
	   .A (new_n11784_) );
   INV_X1 g5054 (
	   .ZN (new_n11785_),
	   .A (_net_5980) );
   INV_X1 g5053 (
	   .ZN (new_n11784_),
	   .A (_net_6048) );
   MUX2_X1 g5052 (
	   .Z (n8840),
	   .S (new_n7544_),
	   .B (_net_7664),
	   .A (new_n7501_1_) );
   CLKBUF_X1 g5051 (
	   .Z (n8835),
	   .A (_net_7811) );
   OAI221_X1 g5050 (
	   .ZN (n8831),
	   .C2 (new_n7306_),
	   .C1 (new_n11456_),
	   .B2 (new_n7302_1_),
	   .B1 (new_n10222_),
	   .A (new_n11780_) );
   AOI22_X1 g5049 (
	   .ZN (new_n11780_),
	   .B2 (_net_7403),
	   .B1 (new_n9203_),
	   .A2 (_net_7435),
	   .A1 (new_n8694_1_) );
   CLKBUF_X1 g5048 (
	   .Z (n8826),
	   .A (_net_7822) );
   CLKBUF_X1 g5047 (
	   .Z (n8823),
	   .A (net_7542) );
   OAI21_X1 g5046 (
	   .ZN (n8818),
	   .B2 (new_n7646_),
	   .B1 (new_n11776_),
	   .A (new_n11775_) );
   INV_X1 g5045 (
	   .ZN (new_n11776_),
	   .A (_net_7409) );
   NAND2_X1 g5044 (
	   .ZN (new_n11775_),
	   .A2 (new_n7276_),
	   .A1 (new_n7645_) );
   CLKBUF_X1 g5043 (
	   .Z (n8813),
	   .A (_net_7797) );
   NAND4_X1 g5042 (
	   .ZN (n8809),
	   .A4 (_net_6414),
	   .A3 (net_6412),
	   .A2 (new_n11535_),
	   .A1 (new_n11772_) );
   INV_X1 g5041 (
	   .ZN (new_n11772_),
	   .A (_net_6415) );
   CLKBUF_X1 g5040 (
	   .Z (n8805),
	   .A (net_6982) );
   CLKBUF_X1 g5039 (
	   .Z (n8800),
	   .A (_net_7808) );
   CLKBUF_X1 g5038 (
	   .Z (n8797),
	   .A (net_6457) );
   CLKBUF_X1 g5037 (
	   .Z (n8793),
	   .A (net_6882) );
   CLKBUF_X1 g5036 (
	   .Z (n8788),
	   .A (_net_7808) );
   CLKBUF_X1 g5035 (
	   .Z (n8784),
	   .A (x1390) );
   OAI21_X1 g5034 (
	   .ZN (n8780),
	   .B2 (new_n6957_1_),
	   .B1 (new_n11764_),
	   .A (new_n11763_) );
   INV_X1 g5033 (
	   .ZN (new_n11764_),
	   .A (_net_7265) );
   NAND2_X1 g5032 (
	   .ZN (new_n11763_),
	   .A2 (new_n9560_),
	   .A1 (new_n6948_) );
   OAI22_X1 g5031 (
	   .ZN (n8775),
	   .B2 (new_n11761_),
	   .B1 (new_n11760_),
	   .A2 (new_n11759_),
	   .A1 (new_n11758_) );
   XNOR2_X1 g5030 (
	   .ZN (new_n11761_),
	   .B (_net_7230),
	   .A (new_n7676_1_) );
   INV_X1 g5029 (
	   .ZN (new_n11760_),
	   .A (new_n8379_) );
   NOR2_X1 g5028 (
	   .ZN (new_n11759_),
	   .A2 (_net_7230),
	   .A1 (new_n7844_) );
   AOI21_X1 g5027 (
	   .ZN (new_n11758_),
	   .B2 (new_n7843_),
	   .B1 (new_n7813_),
	   .A (new_n11757_) );
   NAND2_X1 g5026 (
	   .ZN (new_n11757_),
	   .A2 (_net_7230),
	   .A1 (new_n7692_) );
   NAND2_X1 g5025 (
	   .ZN (n8771),
	   .A2 (new_n8183_1_),
	   .A1 (new_n11755_) );
   OAI211_X1 g5024 (
	   .ZN (new_n11755_),
	   .C2 (_net_6408),
	   .C1 (new_n9684_),
	   .B (_net_6409),
	   .A (_net_6410) );
   CLKBUF_X1 g5023 (
	   .Z (n8767),
	   .A (net_7110) );
   AND2_X1 g5022 (
	   .ZN (n8762),
	   .A2 (_net_6288),
	   .A1 (new_n7235_1_) );
   CLKBUF_X1 g5021 (
	   .Z (n8757),
	   .A (net_140) );
   MUX2_X1 g5020 (
	   .Z (n8753),
	   .S (new_n7028_),
	   .B (_net_7585),
	   .A (new_n8336_) );
   OAI21_X1 g5019 (
	   .ZN (n8748),
	   .B2 (new_n6897_),
	   .B1 (new_n7527_1_),
	   .A (new_n11749_) );
   NAND2_X1 g5018 (
	   .ZN (new_n11749_),
	   .A2 (new_n7649_1_),
	   .A1 (new_n6896_) );
   MUX2_X1 g5017 (
	   .Z (n8743),
	   .S (new_n6823_),
	   .B (_net_6043),
	   .A (_net_7805) );
   CLKBUF_X1 g5016 (
	   .Z (n8739),
	   .A (net_7389) );
   AND2_X1 g5015 (
	   .ZN (n8734),
	   .A2 (net_340),
	   .A1 (new_n7102_1_) );
   NAND4_X1 g5014 (
	   .ZN (n8730),
	   .A4 (new_n11744_),
	   .A3 (new_n11743_),
	   .A2 (new_n11742_),
	   .A1 (new_n11741_) );
   NAND2_X1 g5013 (
	   .ZN (new_n11744_),
	   .A2 (new_n8738_),
	   .A1 (new_n7556_) );
   AOI22_X1 g5012 (
	   .ZN (new_n11743_),
	   .B2 (_net_6109),
	   .B1 (new_n7210_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n10824_) );
   NAND2_X1 g5011 (
	   .ZN (new_n11742_),
	   .A2 (new_n7565_),
	   .A1 (new_n8275_) );
   NAND2_X1 g5010 (
	   .ZN (new_n11741_),
	   .A2 (new_n7587_),
	   .A1 (new_n8271_1_) );
   OAI211_X1 g5009 (
	   .ZN (n8725),
	   .C2 (new_n7211_),
	   .C1 (new_n7568_),
	   .B (new_n11739_),
	   .A (new_n11738_) );
   NAND3_X1 g5008 (
	   .ZN (new_n11739_),
	   .A3 (new_n9632_),
	   .A2 (new_n9627_),
	   .A1 (new_n7560_) );
   OAI21_X1 g5007 (
	   .ZN (new_n11738_),
	   .B2 (new_n7191_),
	   .B1 (new_n7194_1_),
	   .A (new_n8765_) );
   OAI21_X1 g5006 (
	   .ZN (n8720),
	   .B2 (new_n6897_),
	   .B1 (new_n10691_),
	   .A (new_n11736_) );
   NAND2_X1 g5005 (
	   .ZN (new_n11736_),
	   .A2 (new_n8679_),
	   .A1 (new_n6896_) );
   CLKBUF_X1 g5004 (
	   .Z (n8715),
	   .A (net_6388) );
   NOR2_X1 g5003 (
	   .ZN (n8711),
	   .A2 (new_n8678_),
	   .A1 (new_n8543_) );
   NAND3_X1 g5002 (
	   .ZN (n8708),
	   .A3 (new_n11732_),
	   .A2 (new_n11731_),
	   .A1 (new_n11723_) );
   OR2_X1 g5001 (
	   .ZN (new_n11732_),
	   .A2 (new_n6978_),
	   .A1 (new_n7365_) );
   NOR3_X1 g5000 (
	   .ZN (new_n11731_),
	   .A3 (new_n11730_),
	   .A2 (new_n11726_),
	   .A1 (new_n11724_) );
   NAND3_X1 g4999 (
	   .ZN (new_n11730_),
	   .A3 (new_n11729_),
	   .A2 (new_n11728_),
	   .A1 (new_n11727_) );
   NAND4_X1 g4998 (
	   .ZN (new_n11729_),
	   .A4 (net_167),
	   .A3 (x1231),
	   .A2 (new_n7394_),
	   .A1 (new_n7392_) );
   NAND3_X1 g4997 (
	   .ZN (new_n11728_),
	   .A3 (net_204),
	   .A2 (new_n7388_),
	   .A1 (new_n7386_1_) );
   NAND3_X1 g4996 (
	   .ZN (new_n11727_),
	   .A3 (net_241),
	   .A2 (new_n7382_),
	   .A1 (new_n7380_) );
   OAI22_X1 g4995 (
	   .ZN (new_n11726_),
	   .B2 (new_n7377_),
	   .B1 (new_n10136_),
	   .A2 (new_n11725_),
	   .A1 (new_n7374_) );
   INV_X1 g4994 (
	   .ZN (new_n11725_),
	   .A (_net_125) );
   AND4_X1 g4993 (
	   .ZN (new_n11724_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7357_),
	   .A1 (_net_6042) );
   NOR2_X1 g4992 (
	   .ZN (new_n11723_),
	   .A2 (new_n11722_),
	   .A1 (new_n11721_) );
   NOR2_X1 g4991 (
	   .ZN (new_n11722_),
	   .A2 (new_n6901_),
	   .A1 (new_n7362_) );
   NOR2_X1 g4990 (
	   .ZN (new_n11721_),
	   .A2 (new_n11720_),
	   .A1 (new_n9215_1_) );
   INV_X1 g4989 (
	   .ZN (new_n11720_),
	   .A (_net_7702) );
   MUX2_X1 g4988 (
	   .Z (n8703),
	   .S (new_n7436_),
	   .B (_net_6010),
	   .A (_net_7813) );
   CLKBUF_X1 g4987 (
	   .Z (n8698),
	   .A (x1451) );
   OAI21_X1 g4986 (
	   .ZN (n8694),
	   .B2 (new_n7292_1_),
	   .B1 (new_n11716_),
	   .A (new_n11715_) );
   INV_X1 g4985 (
	   .ZN (new_n11716_),
	   .A (_net_6144) );
   NAND2_X1 g4984 (
	   .ZN (new_n11715_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n9746_1_) );
   MUX2_X1 g4983 (
	   .Z (n8689),
	   .S (new_n7503_),
	   .B (_net_7627),
	   .A (new_n7022_) );
   CLKBUF_X1 g4982 (
	   .Z (n8685),
	   .A (net_6722) );
   CLKBUF_X1 g4981 (
	   .Z (n8681),
	   .A (net_6891) );
   NOR2_X1 g4980 (
	   .ZN (n8676),
	   .A2 (_net_6401),
	   .A1 (new_n9442_) );
   OAI21_X1 g4979 (
	   .ZN (n8671),
	   .B2 (new_n6957_1_),
	   .B1 (new_n11709_),
	   .A (new_n11708_) );
   INV_X1 g4978 (
	   .ZN (new_n11709_),
	   .A (_net_7267) );
   NAND2_X1 g4977 (
	   .ZN (new_n11708_),
	   .A2 (new_n7667_),
	   .A1 (new_n6948_) );
   NOR2_X1 g4976 (
	   .ZN (n8666),
	   .A2 (new_n8104_),
	   .A1 (new_n8675_) );
   OAI221_X1 g4975 (
	   .ZN (n8662),
	   .C2 (new_n7306_),
	   .C1 (new_n10266_),
	   .B2 (new_n7302_1_),
	   .B1 (new_n8997_),
	   .A (new_n11705_) );
   AOI22_X1 g4974 (
	   .ZN (new_n11705_),
	   .B2 (_net_7406),
	   .B1 (new_n9203_),
	   .A2 (_net_7438),
	   .A1 (new_n8694_1_) );
   CLKBUF_X1 g4973 (
	   .Z (n8658),
	   .A (net_6600) );
   CLKBUF_X1 g4972 (
	   .Z (n8654),
	   .A (net_6577) );
   CLKBUF_X1 g4971 (
	   .Z (n8650),
	   .A (net_6865) );
   NAND3_X1 g4970 (
	   .ZN (n8645),
	   .A3 (new_n11700_),
	   .A2 (new_n11699_),
	   .A1 (new_n11695_) );
   AOI22_X1 g4969 (
	   .ZN (new_n11700_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6954),
	   .A2 (new_n8457_),
	   .A1 (new_n6879_) );
   AND3_X1 g4968 (
	   .ZN (new_n11699_),
	   .A3 (new_n11698_),
	   .A2 (new_n11697_),
	   .A1 (new_n11696_) );
   NAND2_X1 g4967 (
	   .ZN (new_n11698_),
	   .A2 (_net_6141),
	   .A1 (new_n6868_) );
   NAND2_X1 g4966 (
	   .ZN (new_n11697_),
	   .A2 (new_n6862_),
	   .A1 (new_n8451_1_) );
   NAND2_X1 g4965 (
	   .ZN (new_n11696_),
	   .A2 (new_n6853_),
	   .A1 (new_n10779_) );
   AND3_X1 g4964 (
	   .ZN (new_n11695_),
	   .A3 (new_n11694_),
	   .A2 (new_n11693_),
	   .A1 (new_n11692_) );
   NAND4_X1 g4963 (
	   .ZN (new_n11694_),
	   .A4 (new_n6841_),
	   .A3 (_net_6957),
	   .A2 (net_6922),
	   .A1 (new_n6829_) );
   NAND4_X1 g4962 (
	   .ZN (new_n11693_),
	   .A4 (new_n6836_1_),
	   .A3 (_net_6957),
	   .A2 (net_6858),
	   .A1 (new_n6838_) );
   NAND4_X1 g4961 (
	   .ZN (new_n11692_),
	   .A4 (new_n6833_),
	   .A3 (_net_6957),
	   .A2 (net_6890),
	   .A1 (new_n6830_) );
   CLKBUF_X1 g4960 (
	   .Z (n8641),
	   .A (net_6756) );
   CLKBUF_X1 g4959 (
	   .Z (n8637),
	   .A (net_6013) );
   CLKBUF_X1 g4958 (
	   .Z (n8632),
	   .A (_net_7821) );
   CLKBUF_X1 g4957 (
	   .Z (n8628),
	   .A (_net_7814) );
   AOI21_X1 g4956 (
	   .ZN (n8625),
	   .B2 (new_n8266_1_),
	   .B1 (new_n11686_),
	   .A (new_n8183_1_) );
   NOR2_X1 g4955 (
	   .ZN (new_n11686_),
	   .A2 (_net_6410),
	   .A1 (new_n8187_) );
   CLKBUF_X1 g4954 (
	   .Z (n8621),
	   .A (net_6831) );
   NOR2_X1 g4953 (
	   .ZN (n8616),
	   .A2 (new_n11683_),
	   .A1 (new_n7239_) );
   INV_X1 g4952 (
	   .ZN (new_n11683_),
	   .A (_net_6164) );
   CLKBUF_X1 g4951 (
	   .Z (n8612),
	   .A (net_6463) );
   OAI221_X1 g4950 (
	   .ZN (n8607),
	   .C2 (new_n7312_1_),
	   .C1 (new_n11680_),
	   .B2 (new_n7986_),
	   .B1 (new_n11679_),
	   .A (new_n11678_) );
   INV_X1 g4949 (
	   .ZN (new_n11680_),
	   .A (net_7307) );
   INV_X1 g4948 (
	   .ZN (new_n11679_),
	   .A (net_7371) );
   AOI22_X1 g4947 (
	   .ZN (new_n11678_),
	   .B2 (_net_7275),
	   .B1 (new_n10556_),
	   .A2 (net_7339),
	   .A1 (new_n10555_) );
   OAI21_X1 g4946 (
	   .ZN (n8602),
	   .B2 (new_n7225_),
	   .B1 (new_n11676_),
	   .A (new_n11675_) );
   INV_X1 g4945 (
	   .ZN (new_n11676_),
	   .A (_net_7319) );
   NAND2_X1 g4944 (
	   .ZN (new_n11675_),
	   .A2 (new_n8133_),
	   .A1 (new_n7221_1_) );
   CLKBUF_X1 g4943 (
	   .Z (n8598),
	   .A (net_6695) );
   MUX2_X1 g4942 (
	   .Z (n8593),
	   .S (new_n7284_1_),
	   .B (_net_7695),
	   .A (_net_7797) );
   NOR2_X1 g4941 (
	   .ZN (n8588),
	   .A2 (x889),
	   .A1 (new_n11671_) );
   NAND2_X1 g4940 (
	   .ZN (new_n11671_),
	   .A2 (_net_273),
	   .A1 (n8197) );
   AND2_X1 g4939 (
	   .ZN (n8583),
	   .A2 (_net_6281),
	   .A1 (new_n7235_1_) );
   CLKBUF_X1 g4938 (
	   .Z (n8578),
	   .A (net_6385) );
   CLKBUF_X1 g4937 (
	   .Z (n8575),
	   .A (net_6475) );
   MUX2_X1 g4936 (
	   .Z (n8570),
	   .S (_net_154),
	   .B (net_318),
	   .A (_net_122) );
   CLKBUF_X1 g4935 (
	   .Z (n8565),
	   .A (_net_7797) );
   CLKBUF_X1 g4934 (
	   .Z (n8561),
	   .A (_net_7824) );
   OAI221_X1 g4933 (
	   .ZN (n8557),
	   .C2 (new_n6920_),
	   .C1 (new_n11663_),
	   .B2 (new_n6917_),
	   .B1 (new_n10133_),
	   .A (new_n11662_) );
   INV_X1 g4932 (
	   .ZN (new_n11663_),
	   .A (_net_7356) );
   AOI22_X1 g4931 (
	   .ZN (new_n11662_),
	   .B2 (_net_7260),
	   .B1 (new_n10556_),
	   .A2 (_net_7324),
	   .A1 (new_n10555_) );
   CLKBUF_X1 g4930 (
	   .Z (n8552),
	   .A (_net_7795) );
   CLKBUF_X1 g4929 (
	   .Z (n8549),
	   .A (net_6707) );
   CLKBUF_X1 g4928 (
	   .Z (n8544),
	   .A (_net_7804) );
   NAND2_X1 g4927 (
	   .ZN (n8540),
	   .A2 (new_n11657_),
	   .A1 (new_n11656_) );
   AOI22_X1 g4926 (
	   .ZN (new_n11657_),
	   .B2 (new_n6751_),
	   .B1 (_net_7561),
	   .A2 (_net_7657),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g4925 (
	   .ZN (new_n11656_),
	   .B2 (_net_7625),
	   .B1 (new_n8009_),
	   .A2 (new_n7350_),
	   .A1 (_net_7593) );
   CLKBUF_X1 g4924 (
	   .Z (n8535),
	   .A (_net_7806) );
   OAI21_X1 g4923 (
	   .ZN (n8531),
	   .B2 (new_n7252_1_),
	   .B1 (new_n11405_),
	   .A (new_n11653_) );
   NAND2_X1 g4922 (
	   .ZN (new_n11653_),
	   .A2 (new_n6954_),
	   .A1 (new_n7251_) );
   OAI21_X1 g4921 (
	   .ZN (n8526),
	   .B2 (new_n7101_),
	   .B1 (new_n10189_),
	   .A (new_n11651_) );
   NAND2_X1 g4920 (
	   .ZN (new_n11651_),
	   .A2 (new_n7255_),
	   .A1 (new_n7100_) );
   CLKBUF_X1 g4919 (
	   .Z (n8522),
	   .A (net_6838) );
   MUX2_X1 g4918 (
	   .Z (n8517),
	   .S (new_n10364_),
	   .B (_net_7575),
	   .A (n793) );
   CLKBUF_X1 g4917 (
	   .Z (n8513),
	   .A (net_6744) );
   NOR3_X1 g4916 (
	   .ZN (n8508),
	   .A3 (new_n6811_),
	   .A2 (new_n11646_),
	   .A1 (new_n10468_) );
   AOI21_X1 g4915 (
	   .ZN (new_n11646_),
	   .B2 (net_6556),
	   .B1 (_net_5963),
	   .A (_net_6557) );
   CLKBUF_X1 g4914 (
	   .Z (n8504),
	   .A (net_6622) );
   MUX2_X1 g4913 (
	   .Z (n8499),
	   .S (new_n6823_),
	   .B (_net_6039),
	   .A (_net_7801) );
   CLKBUF_X1 g4912 (
	   .Z (n8494),
	   .A (_net_7810) );
   CLKBUF_X1 g4911 (
	   .Z (n8491),
	   .A (net_7020) );
   NAND3_X1 g4910 (
	   .ZN (n8486),
	   .A3 (new_n11640_),
	   .A2 (new_n11634_),
	   .A1 (new_n11630_) );
   AOI22_X1 g4909 (
	   .ZN (new_n11640_),
	   .B2 (net_7221),
	   .B1 (new_n7844_),
	   .A2 (new_n11639_),
	   .A1 (new_n7837_) );
   NAND4_X1 g4908 (
	   .ZN (new_n11639_),
	   .A4 (new_n11638_),
	   .A3 (new_n11637_),
	   .A2 (new_n11636_),
	   .A1 (new_n11635_) );
   NAND3_X1 g4907 (
	   .ZN (new_n11638_),
	   .A3 (net_7205),
	   .A2 (_net_7228),
	   .A1 (_net_7229) );
   NAND3_X1 g4906 (
	   .ZN (new_n11637_),
	   .A3 (net_7173),
	   .A2 (_net_7229),
	   .A1 (new_n7823_) );
   NAND3_X1 g4905 (
	   .ZN (new_n11636_),
	   .A3 (net_7141),
	   .A2 (_net_7228),
	   .A1 (new_n7821_) );
   NAND2_X1 g4904 (
	   .ZN (new_n11635_),
	   .A2 (net_7109),
	   .A1 (new_n7819_) );
   AND3_X1 g4903 (
	   .ZN (new_n11634_),
	   .A3 (new_n11633_),
	   .A2 (new_n11632_),
	   .A1 (new_n11631_) );
   NAND2_X1 g4902 (
	   .ZN (new_n11633_),
	   .A2 (_net_6178),
	   .A1 (new_n7694_) );
   NAND2_X1 g4901 (
	   .ZN (new_n11632_),
	   .A2 (new_n7701_),
	   .A1 (new_n8060_) );
   NAND2_X1 g4900 (
	   .ZN (new_n11631_),
	   .A2 (new_n7690_),
	   .A1 (new_n7842_) );
   AND3_X1 g4899 (
	   .ZN (new_n11630_),
	   .A3 (new_n11629_),
	   .A2 (new_n11628_),
	   .A1 (new_n11627_) );
   NAND4_X1 g4898 (
	   .ZN (new_n11629_),
	   .A4 (new_n7678_),
	   .A3 (net_7189),
	   .A2 (_net_7227),
	   .A1 (new_n7812_) );
   NAND4_X1 g4897 (
	   .ZN (new_n11628_),
	   .A4 (new_n7683_),
	   .A3 (net_7125),
	   .A2 (_net_7227),
	   .A1 (new_n7816_) );
   NAND4_X1 g4896 (
	   .ZN (new_n11627_),
	   .A4 (new_n7681_1_),
	   .A3 (_net_7227),
	   .A2 (net_7157),
	   .A1 (new_n7813_) );
   OAI21_X1 g4895 (
	   .ZN (n8481),
	   .B2 (new_n7272_),
	   .B1 (new_n11625_),
	   .A (new_n11624_) );
   INV_X1 g4894 (
	   .ZN (new_n11625_),
	   .A (_net_7450) );
   NAND2_X1 g4893 (
	   .ZN (new_n11624_),
	   .A2 (new_n9502_1_),
	   .A1 (new_n7271_) );
   CLKBUF_X1 g4892 (
	   .Z (n8477),
	   .A (net_6754) );
   CLKBUF_X1 g4891 (
	   .Z (n8467),
	   .A (_net_7804) );
   CLKBUF_X1 g4890 (
	   .Z (n8464),
	   .A (net_6742) );
   CLKBUF_X1 g4889 (
	   .Z (n8459),
	   .A (_net_7823) );
   CLKBUF_X1 g4888 (
	   .Z (n8455),
	   .A (_net_7813) );
   NOR2_X1 g4887 (
	   .ZN (n8451),
	   .A2 (new_n7594_),
	   .A1 (new_n8543_) );
   AND2_X1 g4886 (
	   .ZN (n8447),
	   .A2 (net_343),
	   .A1 (new_n7102_1_) );
   NOR3_X1 g4885 (
	   .ZN (n8443),
	   .A3 (_net_7688),
	   .A2 (x1155),
	   .A1 (new_n7184_) );
   CLKBUF_X1 g4884 (
	   .Z (n8438),
	   .A (net_391) );
   NAND4_X1 g4883 (
	   .ZN (n8435),
	   .A4 (new_n11613_),
	   .A3 (new_n11612_),
	   .A2 (new_n11611_),
	   .A1 (new_n11610_) );
   NAND4_X1 g4882 (
	   .ZN (new_n11613_),
	   .A4 (net_7712),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7399_) );
   OR2_X1 g4881 (
	   .ZN (new_n11612_),
	   .A2 (new_n7340_1_),
	   .A1 (new_n7365_) );
   OR2_X1 g4880 (
	   .ZN (new_n11611_),
	   .A2 (new_n10244_),
	   .A1 (new_n7361_) );
   NOR2_X1 g4879 (
	   .ZN (new_n11610_),
	   .A2 (new_n11609_),
	   .A1 (new_n11608_) );
   AND2_X1 g4878 (
	   .ZN (new_n11609_),
	   .A2 (net_7741),
	   .A1 (new_n7934_) );
   NAND4_X1 g4877 (
	   .ZN (new_n11608_),
	   .A4 (new_n11607_),
	   .A3 (new_n11606_),
	   .A2 (new_n11605_),
	   .A1 (new_n11604_) );
   NAND4_X1 g4876 (
	   .ZN (new_n11607_),
	   .A4 (_net_177),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g4875 (
	   .ZN (new_n11606_),
	   .A3 (_net_214),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g4874 (
	   .ZN (new_n11605_),
	   .A3 (net_251),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   NAND4_X1 g4873 (
	   .ZN (new_n11604_),
	   .A4 (new_n7354_1_),
	   .A3 (net_151),
	   .A2 (x1261),
	   .A1 (new_n7370_) );
   CLKBUF_X1 g4872 (
	   .Z (n8430),
	   .A (net_6387) );
   NAND4_X1 g4871 (
	   .ZN (n8426),
	   .A4 (new_n11601_),
	   .A3 (new_n11600_),
	   .A2 (new_n11599_),
	   .A1 (new_n11598_) );
   NAND2_X1 g4870 (
	   .ZN (new_n11601_),
	   .A2 (new_n7013_1_),
	   .A1 (new_n8123_) );
   NAND2_X1 g4869 (
	   .ZN (new_n11600_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n8119_) );
   NAND2_X1 g4868 (
	   .ZN (new_n11599_),
	   .A2 (new_n10655_),
	   .A1 (new_n7000_1_) );
   AOI22_X1 g4867 (
	   .ZN (new_n11598_),
	   .B2 (new_n6985_),
	   .B1 (_net_6089),
	   .A2 (new_n6980_),
	   .A1 (new_n11249_) );
   CLKBUF_X1 g4866 (
	   .Z (n8422),
	   .A (net_7237) );
   CLKBUF_X1 g4865 (
	   .Z (n8418),
	   .A (net_6392) );
   CLKBUF_X1 g4864 (
	   .Z (n8415),
	   .A (net_7137) );
   OAI21_X1 g4863 (
	   .ZN (n8410),
	   .B2 (new_n7225_),
	   .B1 (new_n11593_),
	   .A (new_n11592_) );
   INV_X1 g4862 (
	   .ZN (new_n11593_),
	   .A (_net_7333) );
   NAND2_X1 g4861 (
	   .ZN (new_n11592_),
	   .A2 (new_n9707_),
	   .A1 (new_n7221_1_) );
   NOR2_X1 g4860 (
	   .ZN (n8405),
	   .A2 (new_n11590_),
	   .A1 (new_n11589_) );
   NOR3_X1 g4859 (
	   .ZN (new_n11590_),
	   .A3 (new_n8404_),
	   .A2 (_net_6958),
	   .A1 (new_n9255_) );
   NOR3_X1 g4858 (
	   .ZN (new_n11589_),
	   .A3 (new_n6869_),
	   .A2 (new_n6848_),
	   .A1 (new_n6879_) );
   CLKBUF_X1 g4857 (
	   .Z (n8401),
	   .A (net_7104) );
   MUX2_X1 g4856 (
	   .Z (n8396),
	   .S (new_n10364_),
	   .B (_net_7568),
	   .A (new_n7501_1_) );
   CLKBUF_X1 g4855 (
	   .Z (n8392),
	   .A (net_6425) );
   OAI21_X1 g4854 (
	   .ZN (n8387),
	   .B2 (new_n11584_),
	   .B1 (new_n11583_),
	   .A (new_n9546_1_) );
   NAND2_X1 g4853 (
	   .ZN (new_n11584_),
	   .A2 (_net_5975),
	   .A1 (n9778) );
   OAI21_X1 g4852 (
	   .ZN (new_n11583_),
	   .B2 (new_n11582_),
	   .B1 (new_n11581_),
	   .A (new_n11344_) );
   NOR2_X1 g4851 (
	   .ZN (new_n11582_),
	   .A2 (_net_6963),
	   .A1 (new_n8400_) );
   NOR2_X1 g4850 (
	   .ZN (new_n11581_),
	   .A2 (_net_6960),
	   .A1 (new_n8600_) );
   MUX2_X1 g4849 (
	   .Z (n8382),
	   .S (new_n7028_),
	   .B (_net_7602),
	   .A (new_n8001_) );
   AOI21_X1 g4848 (
	   .ZN (n8377),
	   .B2 (new_n11578_),
	   .B1 (new_n7404_1_),
	   .A (new_n7427_1_) );
   INV_X1 g4847 (
	   .ZN (new_n11578_),
	   .A (_net_7735) );
   OAI221_X1 g4846 (
	   .ZN (n8372),
	   .C2 (new_n11576_),
	   .C1 (new_n8327_),
	   .B2 (new_n10093_),
	   .B1 (new_n7027_1_),
	   .A (new_n11574_) );
   NAND2_X1 g4845 (
	   .ZN (new_n11576_),
	   .A2 (new_n10094_1_),
	   .A1 (new_n11575_) );
   OAI21_X1 g4844 (
	   .ZN (new_n11575_),
	   .B2 (new_n7502_),
	   .B1 (new_n7025_),
	   .A (new_n7027_1_) );
   NAND3_X1 g4843 (
	   .ZN (new_n11574_),
	   .A3 (new_n7020_),
	   .A2 (new_n8326_),
	   .A1 (new_n11573_) );
   XOR2_X1 g4842 (
	   .Z (new_n11573_),
	   .B (_net_7685),
	   .A (_net_7684) );
   NOR2_X1 g4841 (
	   .ZN (n8367),
	   .A2 (new_n9464_),
	   .A1 (new_n9463_) );
   AND2_X1 g4840 (
	   .ZN (n8362),
	   .A2 (net_375),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g4839 (
	   .Z (n8359),
	   .A (net_6427) );
   NOR2_X1 g4838 (
	   .ZN (n8354),
	   .A2 (new_n11568_),
	   .A1 (new_n11567_) );
   NOR3_X1 g4837 (
	   .ZN (new_n11568_),
	   .A3 (new_n7570_),
	   .A2 (new_n7210_),
	   .A1 (new_n7565_) );
   NOR3_X1 g4836 (
	   .ZN (new_n11567_),
	   .A3 (_net_6823),
	   .A2 (new_n8765_),
	   .A1 (new_n7556_) );
   CLKBUF_X1 g4835 (
	   .Z (n8350),
	   .A (net_7023) );
   NAND2_X1 g4834 (
	   .ZN (n8345),
	   .A2 (new_n11564_),
	   .A1 (new_n11554_) );
   AND4_X1 g4833 (
	   .ZN (new_n11564_),
	   .A4 (new_n11563_),
	   .A3 (new_n11562_),
	   .A2 (new_n11556_),
	   .A1 (new_n11555_) );
   NAND2_X1 g4832 (
	   .ZN (new_n11563_),
	   .A2 (_net_6123),
	   .A1 (new_n7209_) );
   NAND2_X1 g4831 (
	   .ZN (new_n11562_),
	   .A2 (new_n7202_),
	   .A1 (new_n11561_) );
   NAND4_X1 g4830 (
	   .ZN (new_n11561_),
	   .A4 (new_n11560_),
	   .A3 (new_n11559_),
	   .A2 (new_n11558_),
	   .A1 (new_n11557_) );
   NAND3_X1 g4829 (
	   .ZN (new_n11560_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6809) );
   NAND3_X1 g4828 (
	   .ZN (new_n11559_),
	   .A3 (_net_6824),
	   .A2 (net_6777),
	   .A1 (new_n7570_) );
   NAND3_X1 g4827 (
	   .ZN (new_n11558_),
	   .A3 (_net_6823),
	   .A2 (net_6745),
	   .A1 (new_n7568_) );
   NAND2_X1 g4826 (
	   .ZN (new_n11557_),
	   .A2 (net_6713),
	   .A1 (new_n7566_) );
   NAND2_X1 g4825 (
	   .ZN (new_n11556_),
	   .A2 (new_n7587_),
	   .A1 (new_n8738_) );
   NAND2_X1 g4824 (
	   .ZN (new_n11555_),
	   .A2 (new_n8744_),
	   .A1 (new_n7564_) );
   AND4_X1 g4823 (
	   .ZN (new_n11554_),
	   .A4 (new_n11553_),
	   .A3 (new_n11552_),
	   .A2 (new_n11551_),
	   .A1 (new_n11550_) );
   NAND4_X1 g4822 (
	   .ZN (new_n11553_),
	   .A4 (new_n7193_),
	   .A3 (net_6757),
	   .A2 (_net_6822),
	   .A1 (new_n7559_) );
   NAND4_X1 g4821 (
	   .ZN (new_n11552_),
	   .A4 (new_n7191_),
	   .A3 (net_6789),
	   .A2 (_net_6822),
	   .A1 (new_n7560_) );
   NAND3_X1 g4820 (
	   .ZN (new_n11551_),
	   .A3 (new_n7189_),
	   .A2 (net_6821),
	   .A1 (new_n7555_) );
   NAND3_X1 g4819 (
	   .ZN (new_n11550_),
	   .A3 (new_n7196_),
	   .A2 (net_6725),
	   .A1 (new_n7555_) );
   CLKBUF_X1 g4818 (
	   .Z (n8340),
	   .A (_net_7812) );
   CLKBUF_X1 g4817 (
	   .Z (n8337),
	   .A (_net_7806) );
   CLKBUF_X1 g4816 (
	   .Z (n8334),
	   .A (net_6851) );
   CLKBUF_X1 g4815 (
	   .Z (n8329),
	   .A (_net_6100) );
   AND2_X1 g4814 (
	   .ZN (n8324),
	   .A2 (_net_6200),
	   .A1 (new_n7235_1_) );
   CLKBUF_X1 g4813 (
	   .Z (n8320),
	   .A (net_7138) );
   CLKBUF_X1 g4812 (
	   .Z (n8316),
	   .A (net_6853) );
   CLKBUF_X1 g4811 (
	   .Z (n8311),
	   .A (_net_7816) );
   CLKBUF_X1 g4810 (
	   .Z (n8307),
	   .A (_net_7811) );
   CLKBUF_X1 g4809 (
	   .Z (n8303),
	   .A (_net_7810) );
   MUX2_X1 g4808 (
	   .Z (n8299),
	   .S (new_n7436_),
	   .B (_net_6020),
	   .A (_net_7820) );
   MUX2_X1 g4807 (
	   .Z (n8294),
	   .S (new_n7544_),
	   .B (_net_7648),
	   .A (new_n8899_1_) );
   CLKBUF_X1 g4806 (
	   .Z (n8289),
	   .A (_net_6125) );
   OAI22_X1 g4805 (
	   .ZN (n8284),
	   .B2 (new_n10340_),
	   .B1 (new_n11535_),
	   .A2 (new_n11534_),
	   .A1 (new_n10325_) );
   INV_X1 g4804 (
	   .ZN (new_n11535_),
	   .A (_net_6413) );
   XNOR2_X1 g4803 (
	   .ZN (new_n11534_),
	   .B (_net_6413),
	   .A (net_6412) );
   CLKBUF_X1 g4802 (
	   .Z (n8280),
	   .A (net_7538) );
   CLKBUF_X1 g4801 (
	   .Z (n8276),
	   .A (net_6615) );
   CLKBUF_X1 g4800 (
	   .Z (n8271),
	   .A (_net_6116) );
   CLKBUF_X1 g4799 (
	   .Z (n8266),
	   .A (net_7799) );
   NOR2_X1 g4798 (
	   .ZN (n8262),
	   .A2 (new_n7214_),
	   .A1 (new_n7020_) );
   OAI221_X1 g4797 (
	   .ZN (n8258),
	   .C2 (new_n7306_),
	   .C1 (new_n10940_),
	   .B2 (new_n7302_1_),
	   .B1 (new_n8068_),
	   .A (new_n11527_) );
   AOI22_X1 g4796 (
	   .ZN (new_n11527_),
	   .B2 (_net_7404),
	   .B1 (new_n9203_),
	   .A2 (_net_7436),
	   .A1 (new_n8694_1_) );
   AOI21_X1 g4795 (
	   .ZN (n8253),
	   .B2 (new_n7739_),
	   .B1 (new_n11525_),
	   .A (new_n11524_) );
   INV_X1 g4794 (
	   .ZN (new_n11525_),
	   .A (_net_7432) );
   NOR2_X1 g4793 (
	   .ZN (new_n11524_),
	   .A2 (n5552),
	   .A1 (new_n7738_) );
   CLKBUF_X1 g4792 (
	   .Z (n8249),
	   .A (net_6388) );
   CLKBUF_X1 g4791 (
	   .Z (n8245),
	   .A (net_7799) );
   CLKBUF_X1 g4790 (
	   .Z (n8241),
	   .A (net_6385) );
   MUX2_X1 g4789 (
	   .Z (n8237),
	   .S (new_n10364_),
	   .B (_net_7580),
	   .A (n5814) );
   CLKBUF_X1 g4788 (
	   .Z (n8232),
	   .A (net_7807) );
   CLKBUF_X1 g4787 (
	   .Z (n8228),
	   .A (_net_7810) );
   INV_X1 g4786 (
	   .ZN (n8224),
	   .A (new_n6865_) );
   CLKBUF_X1 g4785 (
	   .Z (n8220),
	   .A (net_6389) );
   MUX2_X1 g4784 (
	   .Z (n8216),
	   .S (new_n7284_1_),
	   .B (_net_7702),
	   .A (_net_7804) );
   AND2_X1 g4783 (
	   .ZN (n8211),
	   .A2 (new_n11513_),
	   .A1 (new_n11512_) );
   INV_X1 g4782 (
	   .ZN (new_n11513_),
	   .A (x1062) );
   AOI211_X1 g4781 (
	   .ZN (new_n11512_),
	   .C2 (new_n7633_),
	   .C1 (new_n7632_),
	   .B (new_n7614_),
	   .A (new_n6811_) );
   CLKBUF_X1 g4780 (
	   .Z (n8206),
	   .A (_net_7816) );
   NAND3_X1 g4779 (
	   .ZN (n8202),
	   .A3 (new_n11509_),
	   .A2 (new_n11508_),
	   .A1 (new_n11504_) );
   AOI22_X1 g4778 (
	   .ZN (new_n11509_),
	   .B2 (new_n8180_),
	   .B1 (net_7087),
	   .A2 (new_n8165_),
	   .A1 (new_n7060_) );
   AND3_X1 g4777 (
	   .ZN (new_n11508_),
	   .A3 (new_n11507_),
	   .A2 (new_n11506_),
	   .A1 (new_n11505_) );
   NAND2_X1 g4776 (
	   .ZN (new_n11507_),
	   .A2 (_net_6159),
	   .A1 (new_n7091_) );
   NAND2_X1 g4775 (
	   .ZN (new_n11506_),
	   .A2 (new_n7069_),
	   .A1 (new_n9972_) );
   NAND2_X1 g4774 (
	   .ZN (new_n11505_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n8535_1_) );
   AND3_X1 g4773 (
	   .ZN (new_n11504_),
	   .A3 (new_n11503_),
	   .A2 (new_n11502_),
	   .A1 (new_n11501_) );
   NAND4_X1 g4772 (
	   .ZN (new_n11503_),
	   .A4 (new_n7044_),
	   .A3 (_net_7092),
	   .A2 (net_7055),
	   .A1 (new_n8154_) );
   NAND4_X1 g4771 (
	   .ZN (new_n11502_),
	   .A4 (new_n7052_),
	   .A3 (_net_7092),
	   .A2 (net_6991),
	   .A1 (new_n8158_) );
   NAND4_X1 g4770 (
	   .ZN (new_n11501_),
	   .A4 (new_n7050_),
	   .A3 (net_7023),
	   .A2 (_net_7092),
	   .A1 (new_n8155_) );
   AOI21_X1 g4769 (
	   .ZN (n8192),
	   .B2 (new_n7326_1_),
	   .B1 (new_n11499_),
	   .A (new_n11498_) );
   INV_X1 g4768 (
	   .ZN (new_n11499_),
	   .A (_net_7275) );
   NOR2_X1 g4767 (
	   .ZN (new_n11498_),
	   .A2 (n2084),
	   .A1 (new_n7325_) );
   CLKBUF_X1 g4766 (
	   .Z (n8188),
	   .A (net_6835) );
   CLKBUF_X1 g4765 (
	   .Z (n8183),
	   .A (net_7802) );
   OAI221_X1 g4764 (
	   .ZN (n8179),
	   .C2 (new_n7312_1_),
	   .C1 (new_n11494_),
	   .B2 (new_n7986_),
	   .B1 (new_n11493_),
	   .A (new_n11492_) );
   INV_X1 g4763 (
	   .ZN (new_n11494_),
	   .A (net_7306) );
   INV_X1 g4762 (
	   .ZN (new_n11493_),
	   .A (net_7370) );
   AOI22_X1 g4761 (
	   .ZN (new_n11492_),
	   .B2 (_net_7274),
	   .B1 (new_n10556_),
	   .A2 (net_7338),
	   .A1 (new_n10555_) );
   CLKBUF_X1 g4760 (
	   .Z (n8174),
	   .A (_net_7820) );
   NAND2_X1 g4759 (
	   .ZN (n8170),
	   .A2 (new_n11489_),
	   .A1 (new_n11488_) );
   AOI22_X1 g4758 (
	   .ZN (new_n11489_),
	   .B2 (net_7525),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7493) );
   AOI22_X1 g4757 (
	   .ZN (new_n11488_),
	   .B2 (_net_7429),
	   .B1 (new_n7298_),
	   .A2 (net_7461),
	   .A1 (new_n7296_) );
   CLKBUF_X1 g4756 (
	   .Z (n8166),
	   .A (net_7715) );
   NAND2_X1 g4755 (
	   .ZN (n8161),
	   .A2 (new_n11485_),
	   .A1 (new_n11484_) );
   AOI22_X1 g4754 (
	   .ZN (new_n11485_),
	   .B2 (new_n6751_),
	   .B1 (_net_7564),
	   .A2 (_net_7660),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g4753 (
	   .ZN (new_n11484_),
	   .B2 (_net_7596),
	   .B1 (new_n7350_),
	   .A2 (new_n6746_1_),
	   .A1 (_net_7628) );
   NOR2_X1 g4752 (
	   .ZN (n8156),
	   .A2 (new_n8103_),
	   .A1 (new_n8675_) );
   NOR2_X1 g4751 (
	   .ZN (n8152),
	   .A2 (new_n8411_),
	   .A1 (new_n11481_) );
   NAND3_X1 g4750 (
	   .ZN (new_n11481_),
	   .A3 (new_n7262_),
	   .A2 (new_n7025_),
	   .A1 (new_n8412_) );
   CLKBUF_X1 g4749 (
	   .Z (n8147),
	   .A (_net_7808) );
   CLKBUF_X1 g4748 (
	   .Z (n8144),
	   .A (net_6571) );
   CLKBUF_X1 g4747 (
	   .Z (n8140),
	   .A (net_7141) );
   MUX2_X1 g4746 (
	   .Z (n8135),
	   .S (new_n7029_),
	   .B (_net_7592),
	   .A (new_n9910_) );
   OAI21_X1 g4745 (
	   .ZN (n8130),
	   .B2 (new_n7258_),
	   .B1 (new_n7987_),
	   .A (new_n11475_) );
   NAND2_X1 g4744 (
	   .ZN (new_n11475_),
	   .A2 (new_n7108_),
	   .A1 (new_n7251_) );
   CLKBUF_X1 g4743 (
	   .Z (n8125),
	   .A (_net_7795) );
   MUX2_X1 g4742 (
	   .Z (n8121),
	   .S (new_n10364_),
	   .B (_net_7562),
	   .A (new_n7806_1_) );
   CLKBUF_X1 g4741 (
	   .Z (n8116),
	   .A (_net_7801) );
   NAND2_X1 g4740 (
	   .ZN (n8112),
	   .A2 (new_n11470_),
	   .A1 (new_n11465_) );
   AND4_X1 g4739 (
	   .ZN (new_n11470_),
	   .A4 (new_n11469_),
	   .A3 (new_n11468_),
	   .A2 (new_n11467_),
	   .A1 (new_n11466_) );
   NAND2_X1 g4738 (
	   .ZN (new_n11469_),
	   .A2 (_net_6115),
	   .A1 (new_n7209_) );
   NAND2_X1 g4737 (
	   .ZN (new_n11468_),
	   .A2 (new_n7586_1_),
	   .A1 (new_n10830_) );
   NAND2_X1 g4736 (
	   .ZN (new_n11467_),
	   .A2 (new_n7202_),
	   .A1 (new_n10741_) );
   NAND2_X1 g4735 (
	   .ZN (new_n11466_),
	   .A2 (new_n10836_),
	   .A1 (new_n7564_) );
   AND4_X1 g4734 (
	   .ZN (new_n11465_),
	   .A4 (new_n11464_),
	   .A3 (new_n11463_),
	   .A2 (new_n11462_),
	   .A1 (new_n11461_) );
   NAND4_X1 g4733 (
	   .ZN (new_n11464_),
	   .A4 (new_n7194_1_),
	   .A3 (net_6749),
	   .A2 (_net_6822),
	   .A1 (new_n7559_) );
   NAND4_X1 g4732 (
	   .ZN (new_n11463_),
	   .A4 (new_n7191_),
	   .A3 (net_6781),
	   .A2 (_net_6822),
	   .A1 (new_n7560_) );
   NAND3_X1 g4731 (
	   .ZN (new_n11462_),
	   .A3 (new_n7189_),
	   .A2 (net_6813),
	   .A1 (new_n7555_) );
   NAND3_X1 g4730 (
	   .ZN (new_n11461_),
	   .A3 (new_n7196_),
	   .A2 (net_6717),
	   .A1 (new_n7556_) );
   OAI21_X1 g4729 (
	   .ZN (n8107),
	   .B2 (new_n7652_),
	   .B1 (new_n11459_),
	   .A (new_n11458_) );
   INV_X1 g4728 (
	   .ZN (new_n11459_),
	   .A (_net_7417) );
   NAND2_X1 g4727 (
	   .ZN (new_n11458_),
	   .A2 (new_n6904_),
	   .A1 (new_n7645_) );
   OAI21_X1 g4726 (
	   .ZN (n8102),
	   .B2 (new_n7736_),
	   .B1 (new_n11456_),
	   .A (new_n11455_) );
   INV_X1 g4725 (
	   .ZN (new_n11456_),
	   .A (_net_7499) );
   NAND2_X1 g4724 (
	   .ZN (new_n11455_),
	   .A2 (new_n9722_),
	   .A1 (new_n7732_1_) );
   MUX2_X1 g4723 (
	   .Z (n8097),
	   .S (new_n10364_),
	   .B (_net_7573),
	   .A (n718) );
   CLKBUF_X1 g4722 (
	   .Z (n8092),
	   .A (_net_7801) );
   CLKBUF_X1 g4721 (
	   .Z (n8088),
	   .A (_net_7808) );
   CLKBUF_X1 g4720 (
	   .Z (n8085),
	   .A (net_6596) );
   OAI21_X1 g4719 (
	   .ZN (n8080),
	   .B2 (new_n6957_1_),
	   .B1 (new_n11449_),
	   .A (new_n11448_) );
   INV_X1 g4718 (
	   .ZN (new_n11449_),
	   .A (_net_7262) );
   NAND2_X1 g4717 (
	   .ZN (new_n11448_),
	   .A2 (new_n8042_1_),
	   .A1 (new_n6948_) );
   CLKBUF_X1 g4716 (
	   .Z (n8075),
	   .A (_net_7824) );
   CLKBUF_X1 g4715 (
	   .Z (n8072),
	   .A (net_6614) );
   CLKBUF_X1 g4714 (
	   .Z (n8067),
	   .A (_net_7813) );
   CLKBUF_X1 g4713 (
	   .Z (n8064),
	   .A (net_6968) );
   CLKBUF_X1 g4712 (
	   .Z (n8059),
	   .A (_net_7819) );
   CLKBUF_X1 g4711 (
	   .Z (n8056),
	   .A (net_6988) );
   CLKBUF_X1 g4710 (
	   .Z (n8051),
	   .A (net_6399) );
   CLKBUF_X1 g4709 (
	   .Z (n8047),
	   .A (_net_6169) );
   NAND2_X1 g4708 (
	   .ZN (n8042),
	   .A2 (n4304),
	   .A1 (new_n7422_1_) );
   NOR2_X1 g4707 (
	   .ZN (n8038),
	   .A2 (new_n8325_),
	   .A1 (new_n6960_1_) );
   NAND3_X1 g4706 (
	   .ZN (n8033),
	   .A3 (new_n11436_),
	   .A2 (new_n11432_),
	   .A1 (new_n11431_) );
   AND3_X1 g4705 (
	   .ZN (new_n11436_),
	   .A3 (new_n11435_),
	   .A2 (new_n11434_),
	   .A1 (new_n11433_) );
   NAND2_X1 g4704 (
	   .ZN (new_n11435_),
	   .A2 (_net_6072),
	   .A1 (new_n6812_) );
   NAND2_X1 g4703 (
	   .ZN (new_n11434_),
	   .A2 (new_n6800_),
	   .A1 (new_n8211_1_) );
   NAND2_X1 g4702 (
	   .ZN (new_n11433_),
	   .A2 (new_n6809_1_),
	   .A1 (new_n10625_) );
   AOI22_X1 g4701 (
	   .ZN (new_n11432_),
	   .B2 (net_6540),
	   .B1 (new_n6779_1_),
	   .A2 (new_n6784_),
	   .A1 (new_n8203_) );
   AND3_X1 g4700 (
	   .ZN (new_n11431_),
	   .A3 (new_n11430_),
	   .A2 (new_n11429_),
	   .A1 (new_n11428_) );
   NAND4_X1 g4699 (
	   .ZN (new_n11430_),
	   .A4 (new_n6775_),
	   .A3 (_net_6552),
	   .A2 (net_6508),
	   .A1 (new_n6763_) );
   NAND4_X1 g4698 (
	   .ZN (new_n11429_),
	   .A4 (new_n6770_1_),
	   .A3 (_net_6552),
	   .A2 (net_6444),
	   .A1 (new_n6772_) );
   NAND4_X1 g4697 (
	   .ZN (new_n11428_),
	   .A4 (new_n6767_),
	   .A3 (_net_6552),
	   .A2 (net_6476),
	   .A1 (new_n6764_) );
   CLKBUF_X1 g4696 (
	   .Z (n8028),
	   .A (_net_7815) );
   AND2_X1 g4695 (
	   .ZN (n8024),
	   .A2 (_net_6286),
	   .A1 (new_n7235_1_) );
   MUX2_X1 g4694 (
	   .Z (n8019),
	   .S (new_n7537_),
	   .B (_net_291),
	   .A (_net_7811) );
   CLKBUF_X1 g4693 (
	   .Z (n8015),
	   .A (net_7131) );
   AOI21_X1 g4692 (
	   .ZN (n8010),
	   .B2 (new_n11422_),
	   .B1 (new_n11421_),
	   .A (x889) );
   INV_X1 g4691 (
	   .ZN (new_n11422_),
	   .A (_net_5852) );
   NAND3_X1 g4690 (
	   .ZN (new_n11421_),
	   .A3 (net_7778),
	   .A2 (_net_273),
	   .A1 (n8197) );
   AOI21_X1 g4689 (
	   .ZN (n8197),
	   .B2 (new_n11419_),
	   .B1 (new_n11418_),
	   .A (new_n8193_) );
   AOI21_X1 g4688 (
	   .ZN (new_n11419_),
	   .B2 (new_n11417_),
	   .B1 (new_n11416_),
	   .A (_net_189) );
   OAI21_X1 g4687 (
	   .ZN (new_n11418_),
	   .B2 (new_n11417_),
	   .B1 (new_n11416_),
	   .A (new_n10792_) );
   INV_X1 g4686 (
	   .ZN (new_n11417_),
	   .A (_net_192) );
   NOR2_X1 g4685 (
	   .ZN (new_n11416_),
	   .A2 (_net_271),
	   .A1 (_net_191) );
   CLKBUF_X1 g4684 (
	   .Z (n8005),
	   .A (net_6394) );
   CLKBUF_X1 g4683 (
	   .Z (n8002),
	   .A (net_6975) );
   CLKBUF_X1 g4682 (
	   .Z (n7997),
	   .A (_net_7820) );
   CLKBUF_X1 g4681 (
	   .Z (n7994),
	   .A (net_6585) );
   CLKBUF_X1 g4680 (
	   .Z (n7989),
	   .A (_net_7821) );
   AOI21_X1 g4679 (
	   .ZN (n7985),
	   .B2 (new_n7739_),
	   .B1 (new_n11409_),
	   .A (new_n11408_) );
   INV_X1 g4678 (
	   .ZN (new_n11409_),
	   .A (_net_7425) );
   NOR2_X1 g4677 (
	   .ZN (new_n11408_),
	   .A2 (n2958),
	   .A1 (new_n7738_) );
   OAI221_X1 g4676 (
	   .ZN (n7980),
	   .C2 (new_n6920_),
	   .C1 (new_n11406_),
	   .B2 (new_n6917_),
	   .B1 (new_n11405_),
	   .A (new_n11404_) );
   INV_X1 g4675 (
	   .ZN (new_n11406_),
	   .A (_net_7348) );
   INV_X1 g4674 (
	   .ZN (new_n11405_),
	   .A (_net_7284) );
   AOI22_X1 g4673 (
	   .ZN (new_n11404_),
	   .B2 (_net_7252),
	   .B1 (new_n10556_),
	   .A2 (_net_7316),
	   .A1 (new_n10555_) );
   NOR2_X1 g4672 (
	   .ZN (n7975),
	   .A2 (x977),
	   .A1 (new_n11402_) );
   AOI21_X1 g4671 (
	   .ZN (new_n11402_),
	   .B2 (net_7775),
	   .B1 (new_n9392_),
	   .A (_net_5855) );
   NOR2_X1 g4670 (
	   .ZN (n7970),
	   .A2 (new_n7594_),
	   .A1 (new_n8543_) );
   CLKBUF_X1 g4669 (
	   .Z (n7967),
	   .A (net_6992) );
   CLKBUF_X1 g4668 (
	   .Z (n7962),
	   .A (_net_7811) );
   CLKBUF_X1 g4667 (
	   .Z (n7958),
	   .A (net_138) );
   CLKBUF_X1 g4666 (
	   .Z (n7955),
	   .A (net_6724) );
   AOI21_X1 g4665 (
	   .ZN (n7950),
	   .B2 (net_304),
	   .B1 (_net_6040),
	   .A (new_n11395_) );
   NAND3_X1 g4664 (
	   .ZN (new_n11395_),
	   .A3 (_net_6039),
	   .A2 (new_n11394_),
	   .A1 (new_n7655_) );
   INV_X1 g4663 (
	   .ZN (new_n11394_),
	   .A (net_7760) );
   CLKBUF_X1 g4662 (
	   .Z (n7945),
	   .A (net_6390) );
   CLKBUF_X1 g4661 (
	   .Z (n7942),
	   .A (net_7540) );
   CLKBUF_X1 g4660 (
	   .Z (n7937),
	   .A (_net_7798) );
   NAND2_X1 g4659 (
	   .ZN (n7933),
	   .A2 (new_n11389_),
	   .A1 (new_n11388_) );
   AOI22_X1 g4658 (
	   .ZN (new_n11389_),
	   .B2 (new_n6751_),
	   .B1 (_net_7559),
	   .A2 (_net_7655),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g4657 (
	   .ZN (new_n11388_),
	   .B2 (_net_7623),
	   .B1 (new_n8009_),
	   .A2 (new_n7350_),
	   .A1 (_net_7591) );
   CLKBUF_X1 g4656 (
	   .Z (n7929),
	   .A (net_6568) );
   NOR2_X1 g4655 (
	   .ZN (n7924),
	   .A2 (new_n6933_),
	   .A1 (new_n8543_) );
   CLKBUF_X1 g4654 (
	   .Z (n7920),
	   .A (net_6386) );
   CLKBUF_X1 g4653 (
	   .Z (n7916),
	   .A (_net_6167) );
   AOI21_X1 g4652 (
	   .ZN (n7911),
	   .B2 (new_n11381_),
	   .B1 (new_n7859_),
	   .A (new_n11382_) );
   OAI21_X1 g4651 (
	   .ZN (new_n11382_),
	   .B2 (new_n7859_),
	   .B1 (new_n11381_),
	   .A (_net_5984) );
   NAND2_X1 g4650 (
	   .ZN (new_n11381_),
	   .A2 (new_n6761_1_),
	   .A1 (new_n6781_) );
   CLKBUF_X1 g4649 (
	   .Z (n7906),
	   .A (_net_7822) );
   MUX2_X1 g4648 (
	   .Z (n7902),
	   .S (new_n6823_),
	   .B (_net_6031),
	   .A (_net_7796) );
   NOR2_X1 g4647 (
	   .ZN (n7897),
	   .A2 (x837),
	   .A1 (new_n11377_) );
   AOI21_X1 g4646 (
	   .ZN (new_n11377_),
	   .B2 (net_7780),
	   .B1 (new_n10249_),
	   .A (_net_5850) );
   CLKBUF_X1 g4645 (
	   .Z (n7893),
	   .A (net_7249) );
   OAI21_X1 g4644 (
	   .ZN (n7888),
	   .B2 (new_n6907_),
	   .B1 (new_n7300_),
	   .A (new_n11374_) );
   NAND2_X1 g4643 (
	   .ZN (new_n11374_),
	   .A2 (new_n9901_),
	   .A1 (new_n6896_) );
   CLKBUF_X1 g4642 (
	   .Z (n7883),
	   .A (_net_6148) );
   AND2_X1 g4641 (
	   .ZN (n7878),
	   .A2 (net_379),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g4640 (
	   .Z (n7875),
	   .A (net_6874) );
   CLKBUF_X1 g4639 (
	   .Z (n7871),
	   .A (_net_7800) );
   CLKBUF_X1 g4638 (
	   .Z (n7867),
	   .A (net_6393) );
   OAI21_X1 g4637 (
	   .ZN (n7863),
	   .B2 (new_n10421_),
	   .B1 (new_n11367_),
	   .A (new_n6963_) );
   NOR2_X1 g4636 (
	   .ZN (new_n11367_),
	   .A2 (_net_6409),
	   .A1 (new_n9307_1_) );
   NOR2_X1 g4635 (
	   .ZN (n7858),
	   .A2 (new_n9928_),
	   .A1 (new_n8386_) );
   OAI221_X1 g4634 (
	   .ZN (n7853),
	   .C2 (new_n7306_),
	   .C1 (new_n11364_),
	   .B2 (new_n7303_),
	   .B1 (new_n8231_),
	   .A (new_n11363_) );
   INV_X1 g4633 (
	   .ZN (new_n11364_),
	   .A (_net_7504) );
   AOI22_X1 g4632 (
	   .ZN (new_n11363_),
	   .B2 (_net_7408),
	   .B1 (new_n9203_),
	   .A2 (_net_7440),
	   .A1 (new_n8694_1_) );
   CLKBUF_X1 g4631 (
	   .Z (n7848),
	   .A (net_6382) );
   OAI211_X1 g4630 (
	   .ZN (n7845),
	   .C2 (new_n7366_),
	   .C1 (new_n6867_1_),
	   .B (new_n11360_),
	   .A (new_n11359_) );
   NAND4_X1 g4629 (
	   .ZN (new_n11360_),
	   .A4 (net_7715),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   NOR3_X1 g4628 (
	   .ZN (new_n11359_),
	   .A3 (new_n11358_),
	   .A2 (new_n11357_),
	   .A1 (new_n11355_) );
   AND3_X1 g4627 (
	   .ZN (new_n11358_),
	   .A3 (new_n7382_),
	   .A2 (net_254),
	   .A1 (new_n7380_) );
   NOR2_X1 g4626 (
	   .ZN (new_n11357_),
	   .A2 (new_n11356_),
	   .A1 (new_n7378_) );
   INV_X1 g4625 (
	   .ZN (new_n11356_),
	   .A (net_7744) );
   OAI22_X1 g4624 (
	   .ZN (new_n11355_),
	   .B2 (new_n11354_),
	   .B1 (new_n7938_),
	   .A2 (new_n11353_),
	   .A1 (new_n7936_) );
   INV_X1 g4623 (
	   .ZN (new_n11354_),
	   .A (_net_180) );
   INV_X1 g4622 (
	   .ZN (new_n11353_),
	   .A (_net_217) );
   CLKBUF_X1 g4621 (
	   .Z (n7840),
	   .A (_net_6135) );
   AOI21_X1 g4620 (
	   .ZN (n7835),
	   .B2 (new_n7326_1_),
	   .B1 (new_n11350_),
	   .A (new_n11349_) );
   INV_X1 g4619 (
	   .ZN (new_n11350_),
	   .A (_net_7276) );
   NOR2_X1 g4618 (
	   .ZN (new_n11349_),
	   .A2 (n1639),
	   .A1 (new_n7325_) );
   CLKBUF_X1 g4617 (
	   .Z (n7831),
	   .A (net_6566) );
   CLKBUF_X1 g4616 (
	   .Z (n7826),
	   .A (_net_7801) );
   XNOR2_X1 g4615 (
	   .ZN (n7822),
	   .B (new_n11345_),
	   .A (new_n11344_) );
   NAND2_X1 g4614 (
	   .ZN (new_n11345_),
	   .A2 (net_6961),
	   .A1 (new_n6848_) );
   XNOR2_X1 g4613 (
	   .ZN (new_n11344_),
	   .B (_net_6959),
	   .A (_net_6962) );
   CLKBUF_X1 g4612 (
	   .Z (n7818),
	   .A (net_6386) );
   CLKBUF_X1 g4611 (
	   .Z (n7815),
	   .A (net_6734) );
   CLKBUF_X1 g4610 (
	   .Z (n7810),
	   .A (_net_7797) );
   CLKBUF_X1 g4609 (
	   .Z (n7806),
	   .A (_net_7815) );
   CLKBUF_X1 g4608 (
	   .Z (n7802),
	   .A (_net_7800) );
   OAI21_X1 g4607 (
	   .ZN (n7798),
	   .B2 (new_n7272_),
	   .B1 (new_n11337_),
	   .A (new_n11336_) );
   INV_X1 g4606 (
	   .ZN (new_n11337_),
	   .A (_net_7442) );
   NAND2_X1 g4605 (
	   .ZN (new_n11336_),
	   .A2 (new_n6935_),
	   .A1 (new_n7271_) );
   OAI21_X1 g4604 (
	   .ZN (n7793),
	   .B2 (new_n11334_),
	   .B1 (new_n11333_),
	   .A (new_n11332_) );
   NAND2_X1 g4603 (
	   .ZN (new_n11334_),
	   .A2 (new_n10389_),
	   .A1 (n4276) );
   NAND2_X1 g4602 (
	   .ZN (new_n11333_),
	   .A2 (_net_5983),
	   .A1 (new_n9155_) );
   INV_X1 g4601 (
	   .ZN (new_n11332_),
	   .A (_net_6049) );
   NAND3_X1 g4600 (
	   .ZN (n7788),
	   .A3 (new_n11330_),
	   .A2 (new_n11329_),
	   .A1 (new_n11325_) );
   AOI22_X1 g4599 (
	   .ZN (new_n11330_),
	   .B2 (new_n7136_),
	   .B1 (net_6676),
	   .A2 (new_n7012_),
	   .A1 (new_n11249_) );
   AND3_X1 g4598 (
	   .ZN (new_n11329_),
	   .A3 (new_n11328_),
	   .A2 (new_n11327_),
	   .A1 (new_n11326_) );
   NAND2_X1 g4597 (
	   .ZN (new_n11328_),
	   .A2 (_net_6093),
	   .A1 (new_n6984_) );
   NAND2_X1 g4596 (
	   .ZN (new_n11327_),
	   .A2 (new_n6994_),
	   .A1 (new_n7924_1_) );
   NAND2_X1 g4595 (
	   .ZN (new_n11326_),
	   .A2 (new_n6979_),
	   .A1 (new_n7916_1_) );
   AND3_X1 g4594 (
	   .ZN (new_n11325_),
	   .A3 (new_n11324_),
	   .A2 (new_n11323_),
	   .A1 (new_n11322_) );
   NAND4_X1 g4593 (
	   .ZN (new_n11324_),
	   .A4 (new_n6987_),
	   .A3 (net_6644),
	   .A2 (_net_6687),
	   .A1 (new_n7114_) );
   NAND4_X1 g4592 (
	   .ZN (new_n11323_),
	   .A4 (new_n6990_1_),
	   .A3 (net_6580),
	   .A2 (_net_6687),
	   .A1 (new_n7118_) );
   NAND4_X1 g4591 (
	   .ZN (new_n11322_),
	   .A4 (new_n6989_),
	   .A3 (_net_6687),
	   .A2 (net_6612),
	   .A1 (new_n7115_) );
   CLKBUF_X1 g4590 (
	   .Z (n7784),
	   .A (net_6710) );
   CLKBUF_X1 g4589 (
	   .Z (n7779),
	   .A (_net_7824) );
   CLKBUF_X1 g4588 (
	   .Z (n7776),
	   .A (net_6396) );
   NAND4_X1 g4587 (
	   .ZN (n7773),
	   .A4 (new_n11317_),
	   .A3 (new_n11316_),
	   .A2 (new_n11315_),
	   .A1 (new_n11314_) );
   NAND4_X1 g4586 (
	   .ZN (new_n11317_),
	   .A4 (_net_7707),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   OR2_X1 g4585 (
	   .ZN (new_n11316_),
	   .A2 (new_n7208_),
	   .A1 (new_n7365_) );
   OR2_X1 g4584 (
	   .ZN (new_n11315_),
	   .A2 (new_n8325_),
	   .A1 (new_n7361_) );
   NOR2_X1 g4583 (
	   .ZN (new_n11314_),
	   .A2 (new_n11313_),
	   .A1 (new_n11312_) );
   NOR2_X1 g4582 (
	   .ZN (new_n11313_),
	   .A2 (new_n10305_),
	   .A1 (new_n7378_) );
   NAND4_X1 g4581 (
	   .ZN (new_n11312_),
	   .A4 (new_n11311_),
	   .A3 (new_n11310_),
	   .A2 (new_n11309_),
	   .A1 (new_n11308_) );
   NAND4_X1 g4580 (
	   .ZN (new_n11311_),
	   .A4 (_net_172),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g4579 (
	   .ZN (new_n11310_),
	   .A3 (_net_209),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g4578 (
	   .ZN (new_n11309_),
	   .A3 (net_246),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   NAND4_X1 g4577 (
	   .ZN (new_n11308_),
	   .A4 (new_n7354_1_),
	   .A3 (net_146),
	   .A2 (x1261),
	   .A1 (new_n7370_) );
   MUX2_X1 g4576 (
	   .Z (n7768),
	   .S (new_n7285_),
	   .B (_net_7699),
	   .A (_net_7801) );
   CLKBUF_X1 g4575 (
	   .Z (n7764),
	   .A (net_7160) );
   CLKBUF_X1 g4574 (
	   .Z (n7760),
	   .A (net_7143) );
   CLKBUF_X1 g4573 (
	   .Z (n7756),
	   .A (net_6441) );
   MUX2_X1 g4572 (
	   .Z (n7751),
	   .S (new_n10364_),
	   .B (_net_7555),
	   .A (new_n9197_) );
   AOI21_X1 g4571 (
	   .ZN (n7746),
	   .B2 (new_n8306_),
	   .B1 (_net_6828),
	   .A (new_n11301_) );
   OAI21_X1 g4570 (
	   .ZN (new_n11301_),
	   .B2 (_net_6828),
	   .B1 (new_n8306_),
	   .A (_net_6006) );
   NOR4_X1 g4569 (
	   .ZN (n7741),
	   .A4 (_net_6404),
	   .A3 (new_n8187_),
	   .A2 (new_n9685_),
	   .A1 (new_n9684_) );
   NAND3_X1 g4568 (
	   .ZN (n7737),
	   .A3 (new_n11298_),
	   .A2 (new_n11297_),
	   .A1 (new_n11289_) );
   NAND4_X1 g4567 (
	   .ZN (new_n11298_),
	   .A4 (_net_7703),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR3_X1 g4566 (
	   .ZN (new_n11297_),
	   .A3 (new_n11296_),
	   .A2 (new_n11292_),
	   .A1 (new_n11290_) );
   NAND3_X1 g4565 (
	   .ZN (new_n11296_),
	   .A3 (new_n11295_),
	   .A2 (new_n11294_),
	   .A1 (new_n11293_) );
   NAND4_X1 g4564 (
	   .ZN (new_n11295_),
	   .A4 (net_168),
	   .A3 (x1231),
	   .A2 (new_n7394_),
	   .A1 (new_n7392_) );
   NAND3_X1 g4563 (
	   .ZN (new_n11294_),
	   .A3 (net_205),
	   .A2 (new_n7388_),
	   .A1 (new_n7386_1_) );
   NAND3_X1 g4562 (
	   .ZN (new_n11293_),
	   .A3 (net_242),
	   .A2 (new_n7382_),
	   .A1 (new_n7380_) );
   OAI22_X1 g4561 (
	   .ZN (new_n11292_),
	   .B2 (new_n7377_),
	   .B1 (new_n7429_),
	   .A2 (new_n11291_),
	   .A1 (new_n7374_) );
   INV_X1 g4560 (
	   .ZN (new_n11291_),
	   .A (_net_126) );
   AND4_X1 g4559 (
	   .ZN (new_n11290_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7369_),
	   .A1 (_net_6043) );
   NOR2_X1 g4558 (
	   .ZN (new_n11289_),
	   .A2 (new_n11288_),
	   .A1 (new_n11286_) );
   NOR2_X1 g4557 (
	   .ZN (new_n11288_),
	   .A2 (new_n11287_),
	   .A1 (new_n7365_) );
   INV_X1 g4556 (
	   .ZN (new_n11287_),
	   .A (_net_5999) );
   NOR2_X1 g4555 (
	   .ZN (new_n11286_),
	   .A2 (new_n11285_),
	   .A1 (new_n7362_) );
   INV_X1 g4554 (
	   .ZN (new_n11285_),
	   .A (_net_282) );
   AND2_X1 g4553 (
	   .ZN (n7732),
	   .A2 (net_363),
	   .A1 (new_n6898_) );
   OAI21_X1 g4552 (
	   .ZN (n7728),
	   .B2 (new_n7258_),
	   .B1 (new_n8790_),
	   .A (new_n11282_) );
   NAND2_X1 g4551 (
	   .ZN (new_n11282_),
	   .A2 (new_n9611_1_),
	   .A1 (new_n7251_) );
   AOI21_X1 g4550 (
	   .ZN (n7723),
	   .B2 (new_n7326_1_),
	   .B1 (new_n11280_),
	   .A (new_n11279_) );
   INV_X1 g4549 (
	   .ZN (new_n11280_),
	   .A (_net_7273) );
   NOR2_X1 g4548 (
	   .ZN (new_n11279_),
	   .A2 (n518),
	   .A1 (new_n7325_) );
   CLKBUF_X1 g4547 (
	   .Z (n7719),
	   .A (net_6837) );
   CLKBUF_X1 g4546 (
	   .Z (n7714),
	   .A (_net_226) );
   AOI21_X1 g4545 (
	   .ZN (n7709),
	   .B2 (new_n8759_),
	   .B1 (new_n8758_),
	   .A (new_n8754_) );
   CLKBUF_X1 g4544 (
	   .Z (n7704),
	   .A (_net_6108) );
   CLKBUF_X1 g4543 (
	   .Z (n7700),
	   .A (net_6748) );
   MUX2_X1 g4542 (
	   .Z (n7695),
	   .S (new_n7436_),
	   .B (_net_5995),
	   .A (_net_7801) );
   NAND2_X1 g4541 (
	   .ZN (n7686),
	   .A2 (new_n11271_),
	   .A1 (new_n11270_) );
   AOI22_X1 g4540 (
	   .ZN (new_n11271_),
	   .B2 (_net_7553),
	   .B1 (new_n6751_),
	   .A2 (_net_7617),
	   .A1 (new_n6746_1_) );
   AOI22_X1 g4539 (
	   .ZN (new_n11270_),
	   .B2 (_net_7585),
	   .B1 (new_n7350_),
	   .A2 (new_n7970_1_),
	   .A1 (_net_7649) );
   MUX2_X1 g4538 (
	   .Z (n7681),
	   .S (_net_154),
	   .B (net_321),
	   .A (_net_125) );
   NAND3_X1 g4537 (
	   .ZN (n7676),
	   .A3 (new_n11267_),
	   .A2 (new_n11266_),
	   .A1 (new_n11262_) );
   AOI22_X1 g4536 (
	   .ZN (new_n11267_),
	   .B2 (new_n7136_),
	   .B1 (net_6686),
	   .A2 (new_n10547_),
	   .A1 (new_n7013_1_) );
   AND3_X1 g4535 (
	   .ZN (new_n11266_),
	   .A3 (new_n11265_),
	   .A2 (new_n11264_),
	   .A1 (new_n11263_) );
   NAND2_X1 g4534 (
	   .ZN (new_n11265_),
	   .A2 (_net_6103),
	   .A1 (new_n6984_) );
   NAND2_X1 g4533 (
	   .ZN (new_n11264_),
	   .A2 (new_n6979_),
	   .A1 (new_n11255_) );
   NAND2_X1 g4532 (
	   .ZN (new_n11263_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n10655_) );
   AND3_X1 g4531 (
	   .ZN (new_n11262_),
	   .A3 (new_n11261_),
	   .A2 (new_n11260_),
	   .A1 (new_n11259_) );
   NAND4_X1 g4530 (
	   .ZN (new_n11261_),
	   .A4 (new_n6987_),
	   .A3 (_net_6687),
	   .A2 (net_6654),
	   .A1 (new_n7114_) );
   NAND4_X1 g4529 (
	   .ZN (new_n11260_),
	   .A4 (new_n6990_1_),
	   .A3 (net_6590),
	   .A2 (_net_6687),
	   .A1 (new_n7118_) );
   NAND4_X1 g4528 (
	   .ZN (new_n11259_),
	   .A4 (new_n6989_),
	   .A3 (net_6622),
	   .A2 (_net_6687),
	   .A1 (new_n7115_) );
   NAND4_X1 g4527 (
	   .ZN (n7671),
	   .A4 (new_n11257_),
	   .A3 (new_n11256_),
	   .A2 (new_n11250_),
	   .A1 (new_n11246_) );
   AOI22_X1 g4526 (
	   .ZN (new_n11257_),
	   .B2 (_net_6091),
	   .B1 (new_n6985_),
	   .A2 (new_n6980_),
	   .A1 (new_n7924_1_) );
   NAND2_X1 g4525 (
	   .ZN (new_n11256_),
	   .A2 (new_n11255_),
	   .A1 (new_n7000_1_) );
   NAND4_X1 g4524 (
	   .ZN (new_n11255_),
	   .A4 (new_n11254_),
	   .A3 (new_n11253_),
	   .A2 (new_n11252_),
	   .A1 (new_n11251_) );
   NAND3_X1 g4523 (
	   .ZN (new_n11254_),
	   .A3 (_net_6689),
	   .A2 (net_6674),
	   .A1 (_net_6688) );
   NAND3_X1 g4522 (
	   .ZN (new_n11253_),
	   .A3 (_net_6689),
	   .A2 (net_6642),
	   .A1 (new_n7004_) );
   NAND3_X1 g4521 (
	   .ZN (new_n11252_),
	   .A3 (net_6610),
	   .A2 (_net_6688),
	   .A1 (new_n7002_) );
   NAND2_X1 g4520 (
	   .ZN (new_n11251_),
	   .A2 (net_6578),
	   .A1 (new_n6973_) );
   NAND2_X1 g4519 (
	   .ZN (new_n11250_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n11249_) );
   NAND2_X1 g4518 (
	   .ZN (new_n11249_),
	   .A2 (new_n11248_),
	   .A1 (new_n11247_) );
   AOI22_X1 g4517 (
	   .ZN (new_n11248_),
	   .B2 (net_6564),
	   .B1 (new_n6973_),
	   .A2 (net_6596),
	   .A1 (new_n6971_) );
   AOI22_X1 g4516 (
	   .ZN (new_n11247_),
	   .B2 (net_6660),
	   .B1 (new_n6968_),
	   .A2 (new_n6966_),
	   .A1 (net_6628) );
   NAND2_X1 g4515 (
	   .ZN (new_n11246_),
	   .A2 (new_n7013_1_),
	   .A1 (new_n8119_) );
   AOI21_X1 g4514 (
	   .ZN (n7666),
	   .B2 (new_n11244_),
	   .B1 (new_n11243_),
	   .A (new_n11242_) );
   NOR2_X1 g4513 (
	   .ZN (new_n11244_),
	   .A2 (_net_7228),
	   .A1 (new_n8379_) );
   INV_X1 g4512 (
	   .ZN (new_n11243_),
	   .A (new_n8026_) );
   NOR3_X1 g4511 (
	   .ZN (new_n11242_),
	   .A3 (new_n7823_),
	   .A2 (new_n7694_),
	   .A1 (new_n7836_) );
   NOR2_X1 g4510 (
	   .ZN (n7661),
	   .A2 (new_n6934_1_),
	   .A1 (new_n8543_) );
   CLKBUF_X1 g4509 (
	   .Z (n7658),
	   .A (net_6467) );
   CLKBUF_X1 g4508 (
	   .Z (n7654),
	   .A (net_7139) );
   AND2_X1 g4507 (
	   .ZN (n7649),
	   .A2 (_net_6298),
	   .A1 (new_n7235_1_) );
   CLKBUF_X1 g4506 (
	   .Z (n7644),
	   .A (net_6396) );
   MUX2_X1 g4505 (
	   .Z (n7640),
	   .S (new_n7436_),
	   .B (_net_5999),
	   .A (_net_7805) );
   AND2_X1 g4504 (
	   .ZN (n7635),
	   .A2 (net_374),
	   .A1 (new_n7747_) );
   OAI21_X1 g4503 (
	   .ZN (n7631),
	   .B2 (new_n7225_),
	   .B1 (new_n11233_),
	   .A (new_n11232_) );
   INV_X1 g4502 (
	   .ZN (new_n11233_),
	   .A (_net_7331) );
   NAND2_X1 g4501 (
	   .ZN (new_n11232_),
	   .A2 (new_n7667_),
	   .A1 (new_n7221_1_) );
   NOR2_X1 g4500 (
	   .ZN (n7626),
	   .A2 (new_n8678_),
	   .A1 (new_n8543_) );
   AND2_X1 g4499 (
	   .ZN (n7622),
	   .A2 (_net_6206),
	   .A1 (new_n7235_1_) );
   CLKBUF_X1 g4498 (
	   .Z (n7618),
	   .A (net_7392) );
   OAI221_X1 g4497 (
	   .ZN (n7613),
	   .C2 (new_n7303_),
	   .C1 (new_n11176_),
	   .B2 (new_n7305_),
	   .B1 (new_n7735_),
	   .A (new_n11227_) );
   AOI22_X1 g4496 (
	   .ZN (new_n11227_),
	   .B2 (_net_7407),
	   .B1 (new_n9203_),
	   .A2 (_net_7439),
	   .A1 (new_n8694_1_) );
   OAI221_X1 g4495 (
	   .ZN (n7608),
	   .C2 (new_n8301_),
	   .C1 (new_n6846_),
	   .B2 (new_n8593_1_),
	   .B1 (new_n6877_),
	   .A (new_n11225_) );
   OAI21_X1 g4494 (
	   .ZN (new_n11225_),
	   .B2 (new_n6841_),
	   .B1 (new_n6833_),
	   .A (new_n8404_) );
   CLKBUF_X1 g4493 (
	   .Z (n7604),
	   .A (net_6716) );
   AND2_X1 g4492 (
	   .ZN (n7599),
	   .A2 (net_363),
	   .A1 (new_n6898_) );
   OAI221_X1 g4491 (
	   .ZN (n7596),
	   .C2 (new_n7936_),
	   .C1 (new_n11221_),
	   .B2 (new_n7366_),
	   .B1 (new_n7794_),
	   .A (new_n11220_) );
   INV_X1 g4490 (
	   .ZN (new_n11221_),
	   .A (net_222) );
   AOI22_X1 g4489 (
	   .ZN (new_n11220_),
	   .B2 (net_185),
	   .B1 (new_n9730_),
	   .A2 (new_n9729_1_),
	   .A1 (net_259) );
   MUX2_X1 g4488 (
	   .Z (n7591),
	   .S (_net_154),
	   .B (net_323),
	   .A (_net_127) );
   MUX2_X1 g4487 (
	   .Z (n7586),
	   .S (new_n6823_),
	   .B (_net_6033),
	   .A (_net_7798) );
   CLKBUF_X1 g4486 (
	   .Z (n7581),
	   .A (_net_7814) );
   CLKBUF_X1 g4485 (
	   .Z (n7577),
	   .A (_net_6123) );
   NAND2_X1 g4484 (
	   .ZN (n7572),
	   .A2 (new_n11214_),
	   .A1 (new_n11213_) );
   NAND2_X1 g4483 (
	   .ZN (new_n11214_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n8298_) );
   AOI22_X1 g4482 (
	   .ZN (new_n11213_),
	   .B2 (new_n6869_),
	   .B1 (_net_6127),
	   .A2 (new_n6854_),
	   .A1 (new_n10783_) );
   CLKBUF_X1 g4481 (
	   .Z (n7567),
	   .A (x1345) );
   OAI21_X1 g4480 (
	   .ZN (n7563),
	   .B2 (new_n7258_),
	   .B1 (new_n10576_),
	   .A (new_n11210_) );
   NAND2_X1 g4479 (
	   .ZN (new_n11210_),
	   .A2 (new_n8852_),
	   .A1 (new_n7251_) );
   AOI21_X1 g4478 (
	   .ZN (n7558),
	   .B2 (new_n11208_),
	   .B1 (new_n11207_),
	   .A (new_n11206_) );
   AOI21_X1 g4477 (
	   .ZN (new_n11208_),
	   .B2 (_net_267),
	   .B1 (new_n9619_),
	   .A (new_n6943_1_) );
   NAND2_X1 g4476 (
	   .ZN (new_n11207_),
	   .A2 (new_n6952_1_),
	   .A1 (new_n11205_) );
   AOI21_X1 g4475 (
	   .ZN (new_n11206_),
	   .B2 (new_n7102_1_),
	   .B1 (new_n11205_),
	   .A (_net_7381) );
   NOR2_X1 g4474 (
	   .ZN (new_n11205_),
	   .A2 (new_n8193_),
	   .A1 (new_n9619_) );
   CLKBUF_X1 g4473 (
	   .Z (n7553),
	   .A (_net_6090) );
   NAND2_X1 g4472 (
	   .ZN (n7548),
	   .A2 (new_n11202_),
	   .A1 (new_n11201_) );
   AOI22_X1 g4471 (
	   .ZN (new_n11202_),
	   .B2 (new_n6751_),
	   .B1 (_net_7565),
	   .A2 (_net_7661),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g4470 (
	   .ZN (new_n11201_),
	   .B2 (_net_7597),
	   .B1 (new_n7350_),
	   .A2 (new_n6746_1_),
	   .A1 (_net_7629) );
   OAI221_X1 g4469 (
	   .ZN (n7543),
	   .C2 (new_n6920_),
	   .C1 (new_n11199_),
	   .B2 (new_n6917_),
	   .B1 (new_n11198_),
	   .A (new_n11197_) );
   INV_X1 g4468 (
	   .ZN (new_n11199_),
	   .A (net_7367) );
   INV_X1 g4467 (
	   .ZN (new_n11198_),
	   .A (net_7303) );
   AOI22_X1 g4466 (
	   .ZN (new_n11197_),
	   .B2 (_net_7271),
	   .B1 (new_n10556_),
	   .A2 (net_7335),
	   .A1 (new_n10555_) );
   NAND3_X1 g4465 (
	   .ZN (n7539),
	   .A3 (new_n11195_),
	   .A2 (new_n11194_),
	   .A1 (new_n11186_) );
   NAND4_X1 g4464 (
	   .ZN (new_n11195_),
	   .A4 (_net_7705),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR3_X1 g4463 (
	   .ZN (new_n11194_),
	   .A3 (new_n11193_),
	   .A2 (new_n11189_),
	   .A1 (new_n11187_) );
   NAND3_X1 g4462 (
	   .ZN (new_n11193_),
	   .A3 (new_n11192_),
	   .A2 (new_n11191_),
	   .A1 (new_n11190_) );
   NAND4_X1 g4461 (
	   .ZN (new_n11192_),
	   .A4 (net_170),
	   .A3 (x1231),
	   .A2 (new_n7394_),
	   .A1 (new_n7392_) );
   NAND3_X1 g4460 (
	   .ZN (new_n11191_),
	   .A3 (net_207),
	   .A2 (new_n7388_),
	   .A1 (new_n7386_1_) );
   NAND3_X1 g4459 (
	   .ZN (new_n11190_),
	   .A3 (net_244),
	   .A2 (new_n7382_),
	   .A1 (new_n7380_) );
   OAI22_X1 g4458 (
	   .ZN (new_n11189_),
	   .B2 (new_n7378_),
	   .B1 (new_n10379_),
	   .A2 (new_n11188_),
	   .A1 (new_n7374_) );
   INV_X1 g4457 (
	   .ZN (new_n11188_),
	   .A (_net_128) );
   AND4_X1 g4456 (
	   .ZN (new_n11187_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7369_),
	   .A1 (_net_6045) );
   NOR2_X1 g4455 (
	   .ZN (new_n11186_),
	   .A2 (new_n11185_),
	   .A1 (new_n11183_) );
   NOR2_X1 g4454 (
	   .ZN (new_n11185_),
	   .A2 (new_n11184_),
	   .A1 (new_n7366_) );
   INV_X1 g4453 (
	   .ZN (new_n11184_),
	   .A (_net_6001) );
   NOR2_X1 g4452 (
	   .ZN (new_n11183_),
	   .A2 (new_n11182_),
	   .A1 (new_n7362_) );
   INV_X1 g4451 (
	   .ZN (new_n11182_),
	   .A (_net_284) );
   CLKBUF_X1 g4450 (
	   .Z (n7535),
	   .A (net_6757) );
   CLKBUF_X1 g4449 (
	   .Z (n7530),
	   .A (_net_7808) );
   CLKBUF_X1 g4448 (
	   .Z (n7527),
	   .A (net_6451) );
   CLKBUF_X1 g4447 (
	   .Z (n7522),
	   .A (_net_7809) );
   OAI21_X1 g4446 (
	   .ZN (n7518),
	   .B2 (new_n6907_),
	   .B1 (new_n11176_),
	   .A (new_n11175_) );
   INV_X1 g4445 (
	   .ZN (new_n11176_),
	   .A (_net_7471) );
   NAND2_X1 g4444 (
	   .ZN (new_n11175_),
	   .A2 (new_n7484_),
	   .A1 (new_n6896_) );
   CLKBUF_X1 g4443 (
	   .Z (n7513),
	   .A (_net_7823) );
   CLKBUF_X1 g4442 (
	   .Z (n7509),
	   .A (_net_7809) );
   CLKBUF_X1 g4441 (
	   .Z (n7505),
	   .A (net_6383) );
   NOR2_X1 g4440 (
	   .ZN (n7501),
	   .A2 (new_n7369_),
	   .A1 (new_n10058_) );
   NAND4_X1 g4439 (
	   .ZN (n7496),
	   .A4 (new_n11169_),
	   .A3 (new_n11168_),
	   .A2 (new_n11167_),
	   .A1 (new_n11166_) );
   NAND2_X1 g4438 (
	   .ZN (new_n11169_),
	   .A2 (new_n6784_),
	   .A1 (new_n9830_) );
   NAND2_X1 g4437 (
	   .ZN (new_n11168_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n8199_) );
   NAND2_X1 g4436 (
	   .ZN (new_n11167_),
	   .A2 (new_n6798_),
	   .A1 (new_n8205_) );
   AOI22_X1 g4435 (
	   .ZN (new_n11166_),
	   .B2 (new_n6813_1_),
	   .B1 (_net_6068),
	   .A2 (new_n7166_),
	   .A1 (new_n8203_) );
   CLKBUF_X1 g4434 (
	   .Z (n7492),
	   .A (net_6726) );
   NOR3_X1 g4433 (
	   .ZN (n7487),
	   .A3 (new_n6867_1_),
	   .A2 (new_n11163_),
	   .A1 (new_n8338_) );
   AOI21_X1 g4432 (
	   .ZN (new_n11163_),
	   .B2 (_net_5975),
	   .B1 (net_6961),
	   .A (_net_6962) );
   CLKBUF_X1 g4431 (
	   .Z (n7482),
	   .A (_net_7810) );
   OAI21_X1 g4430 (
	   .ZN (n7478),
	   .B2 (new_n7111_1_),
	   .B1 (new_n11046_),
	   .A (new_n11160_) );
   NAND2_X1 g4429 (
	   .ZN (new_n11160_),
	   .A2 (new_n8133_),
	   .A1 (new_n7100_) );
   AND2_X1 g4428 (
	   .ZN (n7473),
	   .A2 (_net_6221),
	   .A1 (new_n7235_1_) );
   CLKBUF_X1 g4427 (
	   .Z (n7468),
	   .A (_net_6141) );
   CLKBUF_X1 g4426 (
	   .Z (n7463),
	   .A (_net_7814) );
   OAI21_X1 g4425 (
	   .ZN (n7459),
	   .B2 (new_n6957_1_),
	   .B1 (new_n11155_),
	   .A (new_n11154_) );
   INV_X1 g4424 (
	   .ZN (new_n11155_),
	   .A (_net_7263) );
   NAND2_X1 g4423 (
	   .ZN (new_n11154_),
	   .A2 (new_n8105_),
	   .A1 (new_n6948_) );
   MUX2_X1 g4422 (
	   .Z (n7454),
	   .S (new_n7436_),
	   .B (_net_6007),
	   .A (_net_7810) );
   CLKBUF_X1 g4421 (
	   .Z (n7450),
	   .A (net_6740) );
   CLKBUF_X1 g4420 (
	   .Z (n7446),
	   .A (net_6696) );
   CLKBUF_X1 g4419 (
	   .Z (n7442),
	   .A (net_6700) );
   NAND4_X1 g4418 (
	   .ZN (n7437),
	   .A4 (new_n11148_),
	   .A3 (new_n11147_),
	   .A2 (new_n11146_),
	   .A1 (new_n11145_) );
   NAND2_X1 g4417 (
	   .ZN (new_n11148_),
	   .A2 (new_n6784_),
	   .A1 (new_n8146_) );
   NAND2_X1 g4416 (
	   .ZN (new_n11147_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n8142_) );
   NAND2_X1 g4415 (
	   .ZN (new_n11146_),
	   .A2 (new_n9089_),
	   .A1 (new_n8205_) );
   AOI22_X1 g4414 (
	   .ZN (new_n11145_),
	   .B2 (new_n6813_1_),
	   .B1 (_net_6069),
	   .A2 (new_n7166_),
	   .A1 (new_n9871_1_) );
   INV_X1 g4413 (
	   .ZN (n7432),
	   .A (new_n7055_) );
   CLKBUF_X1 g4412 (
	   .Z (n7427),
	   .A (_net_6149) );
   AOI21_X1 g4411 (
	   .ZN (n7422),
	   .B2 (new_n11140_),
	   .B1 (new_n8591_),
	   .A (new_n11141_) );
   OAI21_X1 g4410 (
	   .ZN (new_n11141_),
	   .B2 (new_n8591_),
	   .B1 (new_n11140_),
	   .A (_net_6017) );
   NAND2_X1 g4409 (
	   .ZN (new_n11140_),
	   .A2 (new_n6827_),
	   .A1 (new_n6866_) );
   CLKBUF_X1 g4408 (
	   .Z (n7417),
	   .A (_net_6081) );
   CLKBUF_X1 g4407 (
	   .Z (n7413),
	   .A (net_6994) );
   CLKBUF_X1 g4406 (
	   .Z (n7408),
	   .A (_net_7819) );
   CLKBUF_X1 g4405 (
	   .Z (n7404),
	   .A (_net_7808) );
   OAI21_X1 g4404 (
	   .ZN (n7400),
	   .B2 (new_n6907_),
	   .B1 (new_n10567_),
	   .A (new_n11134_) );
   NAND2_X1 g4403 (
	   .ZN (new_n11134_),
	   .A2 (new_n7276_),
	   .A1 (new_n6896_) );
   MUX2_X1 g4402 (
	   .Z (n7395),
	   .S (_net_154),
	   .B (net_313),
	   .A (_net_117) );
   CLKBUF_X1 g4401 (
	   .Z (n7391),
	   .A (net_7118) );
   OAI21_X1 g4400 (
	   .ZN (n7386),
	   .B2 (new_n7211_),
	   .B1 (new_n11130_),
	   .A (new_n11129_) );
   INV_X1 g4399 (
	   .ZN (new_n11130_),
	   .A (_net_6105) );
   NAND2_X1 g4398 (
	   .ZN (new_n11129_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n8275_) );
   MUX2_X1 g4397 (
	   .Z (n7381),
	   .S (new_n7545_),
	   .B (_net_7666),
	   .A (new_n8001_) );
   CLKBUF_X1 g4396 (
	   .Z (n7376),
	   .A (net_134) );
   CLKBUF_X1 g4395 (
	   .Z (n7372),
	   .A (_net_7798) );
   CLKBUF_X1 g4394 (
	   .Z (n7368),
	   .A (_net_6121) );
   OAI221_X1 g4393 (
	   .ZN (n7363),
	   .C2 (new_n6920_),
	   .C1 (new_n11123_),
	   .B2 (new_n6917_),
	   .B1 (new_n11122_),
	   .A (new_n11121_) );
   INV_X1 g4392 (
	   .ZN (new_n11123_),
	   .A (net_7375) );
   INV_X1 g4391 (
	   .ZN (new_n11122_),
	   .A (net_7311) );
   AOI22_X1 g4390 (
	   .ZN (new_n11121_),
	   .B2 (_net_7279),
	   .B1 (new_n10556_),
	   .A2 (net_7343),
	   .A1 (new_n10555_) );
   CLKBUF_X1 g4389 (
	   .Z (n7359),
	   .A (net_7008) );
   NAND2_X1 g4388 (
	   .ZN (n7354),
	   .A2 (new_n11118_),
	   .A1 (new_n11117_) );
   AOI22_X1 g4387 (
	   .ZN (new_n11118_),
	   .B2 (_net_7572),
	   .B1 (new_n6755_),
	   .A2 (net_7604),
	   .A1 (new_n6743_) );
   AOI22_X1 g4386 (
	   .ZN (new_n11117_),
	   .B2 (net_7636),
	   .B1 (new_n8009_),
	   .A2 (new_n7970_1_),
	   .A1 (net_7668) );
   CLKBUF_X1 g4385 (
	   .Z (n7349),
	   .A (net_6058) );
   CLKBUF_X1 g4384 (
	   .Z (n7344),
	   .A (_net_7803) );
   NAND3_X1 g4383 (
	   .ZN (n7340),
	   .A3 (new_n11113_),
	   .A2 (new_n11112_),
	   .A1 (new_n11108_) );
   AOI22_X1 g4382 (
	   .ZN (new_n11113_),
	   .B2 (net_7222),
	   .B1 (new_n7844_),
	   .A2 (new_n8368_),
	   .A1 (new_n7837_) );
   AND3_X1 g4381 (
	   .ZN (new_n11112_),
	   .A3 (new_n11111_),
	   .A2 (new_n11110_),
	   .A1 (new_n11109_) );
   NAND2_X1 g4380 (
	   .ZN (new_n11111_),
	   .A2 (_net_6179),
	   .A1 (new_n7694_) );
   NAND2_X1 g4379 (
	   .ZN (new_n11110_),
	   .A2 (new_n7701_),
	   .A1 (new_n8362_1_) );
   NAND2_X1 g4378 (
	   .ZN (new_n11109_),
	   .A2 (new_n7690_),
	   .A1 (new_n10495_) );
   AND3_X1 g4377 (
	   .ZN (new_n11108_),
	   .A3 (new_n11107_),
	   .A2 (new_n11106_),
	   .A1 (new_n11105_) );
   NAND4_X1 g4376 (
	   .ZN (new_n11107_),
	   .A4 (new_n7678_),
	   .A3 (net_7190),
	   .A2 (_net_7227),
	   .A1 (new_n7812_) );
   NAND4_X1 g4375 (
	   .ZN (new_n11106_),
	   .A4 (new_n7683_),
	   .A3 (_net_7227),
	   .A2 (net_7126),
	   .A1 (new_n7816_) );
   NAND4_X1 g4374 (
	   .ZN (new_n11105_),
	   .A4 (new_n7681_1_),
	   .A3 (_net_7227),
	   .A2 (net_7158),
	   .A1 (new_n7813_) );
   CLKBUF_X1 g4373 (
	   .Z (n7335),
	   .A (net_5860) );
   CLKBUF_X1 g4372 (
	   .Z (n7330),
	   .A (_net_6088) );
   CLKBUF_X1 g4371 (
	   .Z (n7326),
	   .A (net_6715) );
   OAI21_X1 g4370 (
	   .ZN (n7321),
	   .B2 (new_n7111_1_),
	   .B1 (new_n6918_),
	   .A (new_n11100_) );
   NAND2_X1 g4369 (
	   .ZN (new_n11100_),
	   .A2 (new_n9707_),
	   .A1 (new_n7100_) );
   CLKBUF_X1 g4368 (
	   .Z (n7316),
	   .A (_net_6178) );
   CLKBUF_X1 g4367 (
	   .Z (n7312),
	   .A (net_6869) );
   MUX2_X1 g4366 (
	   .Z (n7307),
	   .S (new_n7285_),
	   .B (_net_7697),
	   .A (net_7799) );
   AND2_X1 g4365 (
	   .ZN (n7302),
	   .A2 (_net_6287),
	   .A1 (new_n9520_1_) );
   MUX2_X1 g4364 (
	   .Z (n7297),
	   .S (new_n6823_),
	   .B (_net_6028),
	   .A (_net_7793) );
   CLKBUF_X1 g4363 (
	   .Z (n7292),
	   .A (x1406) );
   CLKBUF_X1 g4362 (
	   .Z (n7288),
	   .A (net_6397) );
   CLKBUF_X1 g4361 (
	   .Z (n7284),
	   .A (_net_7816) );
   NAND2_X1 g4360 (
	   .ZN (n7280),
	   .A2 (new_n7430_),
	   .A1 (new_n11090_) );
   NAND2_X1 g4359 (
	   .ZN (new_n11090_),
	   .A2 (_net_5972),
	   .A1 (new_n6866_) );
   AND2_X1 g4358 (
	   .ZN (n7275),
	   .A2 (_net_6290),
	   .A1 (new_n9520_1_) );
   NAND4_X1 g4357 (
	   .ZN (n7270),
	   .A4 (new_n11087_),
	   .A3 (new_n11086_),
	   .A2 (new_n11085_),
	   .A1 (new_n11084_) );
   AOI22_X1 g4356 (
	   .ZN (new_n11087_),
	   .B2 (_net_6151),
	   .B1 (new_n7092_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n8179_1_) );
   NAND2_X1 g4355 (
	   .ZN (new_n11086_),
	   .A2 (new_n8527_),
	   .A1 (new_n7073_) );
   NAND2_X1 g4354 (
	   .ZN (new_n11085_),
	   .A2 (new_n7070_),
	   .A1 (new_n10526_) );
   NAND2_X1 g4353 (
	   .ZN (new_n11084_),
	   .A2 (new_n7060_),
	   .A1 (new_n7413_1_) );
   CLKBUF_X1 g4352 (
	   .Z (n7260),
	   .A (_net_7797) );
   CLKBUF_X1 g4351 (
	   .Z (n7256),
	   .A (net_7792) );
   CLKBUF_X1 g4350 (
	   .Z (n7252),
	   .A (_net_7804) );
   CLKBUF_X1 g4349 (
	   .Z (n7249),
	   .A (x1486) );
   OAI22_X1 g4348 (
	   .ZN (n7245),
	   .B2 (new_n11077_),
	   .B1 (new_n9678_1_),
	   .A2 (new_n11076_),
	   .A1 (new_n9679_) );
   NAND2_X1 g4347 (
	   .ZN (new_n11077_),
	   .A2 (new_n11076_),
	   .A1 (new_n9440_) );
   INV_X1 g4346 (
	   .ZN (new_n11076_),
	   .A (_net_6423) );
   OAI21_X1 g4345 (
	   .ZN (n7240),
	   .B2 (new_n7292_1_),
	   .B1 (new_n11074_),
	   .A (new_n11073_) );
   INV_X1 g4344 (
	   .ZN (new_n11074_),
	   .A (_net_6145) );
   NAND2_X1 g4343 (
	   .ZN (new_n11073_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n7417_1_) );
   AND2_X1 g4342 (
	   .ZN (n7235),
	   .A2 (_net_6294),
	   .A1 (new_n9520_1_) );
   CLKBUF_X1 g4341 (
	   .Z (n7230),
	   .A (_net_7823) );
   AND2_X1 g4340 (
	   .ZN (n7226),
	   .A2 (_net_6239),
	   .A1 (new_n9520_1_) );
   AND2_X1 g4339 (
	   .ZN (n7221),
	   .A2 (_net_6210),
	   .A1 (new_n9520_1_) );
   OAI21_X1 g4338 (
	   .ZN (n7216),
	   .B2 (new_n7111_1_),
	   .B1 (new_n7467_),
	   .A (new_n11067_) );
   NAND2_X1 g4337 (
	   .ZN (new_n11067_),
	   .A2 (new_n9560_),
	   .A1 (new_n7100_) );
   CLKBUF_X1 g4336 (
	   .Z (n7212),
	   .A (net_6559) );
   NAND3_X1 g4335 (
	   .ZN (n7207),
	   .A3 (new_n11064_),
	   .A2 (new_n11060_),
	   .A1 (new_n11059_) );
   AND3_X1 g4334 (
	   .ZN (new_n11064_),
	   .A3 (new_n11063_),
	   .A2 (new_n11062_),
	   .A1 (new_n11061_) );
   NAND2_X1 g4333 (
	   .ZN (new_n11063_),
	   .A2 (_net_6080),
	   .A1 (new_n6812_) );
   NAND2_X1 g4332 (
	   .ZN (new_n11062_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n6792_) );
   NAND2_X1 g4331 (
	   .ZN (new_n11061_),
	   .A2 (new_n7166_),
	   .A1 (new_n6798_) );
   AOI22_X1 g4330 (
	   .ZN (new_n11060_),
	   .B2 (new_n9282_1_),
	   .B1 (new_n6784_),
	   .A2 (new_n6779_1_),
	   .A1 (net_6548) );
   AND3_X1 g4329 (
	   .ZN (new_n11059_),
	   .A3 (new_n11058_),
	   .A2 (new_n11057_),
	   .A1 (new_n11056_) );
   NAND4_X1 g4328 (
	   .ZN (new_n11058_),
	   .A4 (new_n6775_),
	   .A3 (_net_6552),
	   .A2 (net_6516),
	   .A1 (new_n6763_) );
   NAND4_X1 g4327 (
	   .ZN (new_n11057_),
	   .A4 (new_n6770_1_),
	   .A3 (_net_6552),
	   .A2 (net_6452),
	   .A1 (new_n6772_) );
   NAND4_X1 g4326 (
	   .ZN (new_n11056_),
	   .A4 (new_n6767_),
	   .A3 (_net_6552),
	   .A2 (net_6484),
	   .A1 (new_n6764_) );
   CLKBUF_X1 g4325 (
	   .Z (n7203),
	   .A (net_6477) );
   CLKBUF_X1 g4324 (
	   .Z (n7199),
	   .A (net_7238) );
   OAI221_X1 g4323 (
	   .ZN (n7194),
	   .C2 (new_n9469_),
	   .C1 (new_n6787_),
	   .B2 (new_n7847_),
	   .B1 (new_n6782_),
	   .A (new_n11052_) );
   OAI21_X1 g4322 (
	   .ZN (new_n11052_),
	   .B2 (new_n6775_),
	   .B1 (new_n6767_),
	   .A (new_n8908_1_) );
   CLKBUF_X1 g4321 (
	   .Z (n7190),
	   .A (net_6430) );
   NOR2_X1 g4320 (
	   .ZN (n7185),
	   .A2 (new_n8103_),
	   .A1 (new_n8675_) );
   CLKBUF_X1 g4319 (
	   .Z (n7182),
	   .A (net_7543) );
   OAI221_X1 g4318 (
	   .ZN (n7177),
	   .C2 (new_n7312_1_),
	   .C1 (new_n11047_),
	   .B2 (new_n7986_),
	   .B1 (new_n11046_),
	   .A (new_n11045_) );
   INV_X1 g4317 (
	   .ZN (new_n11047_),
	   .A (_net_7287) );
   INV_X1 g4316 (
	   .ZN (new_n11046_),
	   .A (_net_7351) );
   AOI22_X1 g4315 (
	   .ZN (new_n11045_),
	   .B2 (_net_7255),
	   .B1 (new_n10556_),
	   .A2 (_net_7319),
	   .A1 (new_n10555_) );
   NOR2_X1 g4314 (
	   .ZN (n7172),
	   .A2 (new_n7878_1_),
	   .A1 (new_n8386_) );
   CLKBUF_X1 g4313 (
	   .Z (n7167),
	   .A (net_141) );
   OAI211_X1 g4312 (
	   .ZN (n7164),
	   .C2 (new_n9215_1_),
	   .C1 (new_n11041_),
	   .B (new_n11040_),
	   .A (new_n11039_) );
   INV_X1 g4311 (
	   .ZN (new_n11041_),
	   .A (_net_7719) );
   NAND4_X1 g4310 (
	   .ZN (new_n11040_),
	   .A4 (new_n7364_),
	   .A3 (_net_6021),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   NOR3_X1 g4309 (
	   .ZN (new_n11039_),
	   .A3 (new_n11038_),
	   .A2 (new_n11037_),
	   .A1 (new_n11036_) );
   AND3_X1 g4308 (
	   .ZN (new_n11038_),
	   .A3 (new_n7382_),
	   .A2 (net_258),
	   .A1 (new_n7380_) );
   NOR2_X1 g4307 (
	   .ZN (new_n11037_),
	   .A2 (new_n8463_),
	   .A1 (new_n7378_) );
   OAI22_X1 g4306 (
	   .ZN (new_n11036_),
	   .B2 (new_n11035_),
	   .B1 (new_n7938_),
	   .A2 (new_n11034_),
	   .A1 (new_n7936_) );
   INV_X1 g4305 (
	   .ZN (new_n11035_),
	   .A (_net_184) );
   INV_X1 g4304 (
	   .ZN (new_n11034_),
	   .A (_net_221) );
   CLKBUF_X1 g4303 (
	   .Z (n7160),
	   .A (net_6862) );
   CLKBUF_X1 g4302 (
	   .Z (n7155),
	   .A (_net_7824) );
   CLKBUF_X1 g4301 (
	   .Z (n7151),
	   .A (_net_7816) );
   CLKBUF_X1 g4300 (
	   .Z (n7147),
	   .A (_net_6073) );
   NOR2_X1 g4299 (
	   .ZN (n7142),
	   .A2 (new_n9900_),
	   .A1 (new_n8543_) );
   AOI21_X1 g4298 (
	   .ZN (n7138),
	   .B2 (new_n11027_),
	   .B1 (new_n11018_),
	   .A (new_n11019_) );
   INV_X1 g4297 (
	   .ZN (new_n11027_),
	   .A (_net_5848) );
   MUX2_X1 g4296 (
	   .Z (n7133),
	   .S (new_n7285_),
	   .B (_net_7705),
	   .A (net_7807) );
   CLKBUF_X1 g4295 (
	   .Z (n7128),
	   .A (_net_7798) );
   CLKBUF_X1 g4294 (
	   .Z (n7125),
	   .A (net_6561) );
   CLKBUF_X1 g4293 (
	   .Z (n7120),
	   .A (_net_7803) );
   CLKBUF_X1 g4292 (
	   .Z (n7116),
	   .A (_net_6133) );
   CLKBUF_X1 g4291 (
	   .Z (n7111),
	   .A (_net_7821) );
   OAI21_X1 g4290 (
	   .ZN (n7107),
	   .B2 (new_n11019_),
	   .B1 (new_n11018_),
	   .A (new_n11017_) );
   INV_X1 g4289 (
	   .ZN (new_n11019_),
	   .A (net_7767) );
   NAND2_X1 g4288 (
	   .ZN (new_n11018_),
	   .A2 (net_7771),
	   .A1 (new_n8911_) );
   NAND2_X1 g4287 (
	   .ZN (new_n11017_),
	   .A2 (net_7769),
	   .A1 (new_n9042_1_) );
   OAI221_X1 g4286 (
	   .ZN (n7102),
	   .C2 (new_n7303_),
	   .C1 (new_n8289_1_),
	   .B2 (new_n7305_),
	   .B1 (new_n7876_),
	   .A (new_n11015_) );
   AOI22_X1 g4285 (
	   .ZN (new_n11015_),
	   .B2 (_net_7401),
	   .B1 (new_n9203_),
	   .A2 (_net_7433),
	   .A1 (new_n8694_1_) );
   CLKBUF_X1 g4284 (
	   .Z (n7098),
	   .A (net_7152) );
   CLKBUF_X1 g4283 (
	   .Z (n7093),
	   .A (net_6398) );
   CLKBUF_X1 g4282 (
	   .Z (n7089),
	   .A (_net_7811) );
   AND2_X1 g4281 (
	   .ZN (n7085),
	   .A2 (net_361),
	   .A1 (new_n6898_) );
   CLKBUF_X1 g4280 (
	   .Z (n7082),
	   .A (net_6872) );
   AND2_X1 g4279 (
	   .ZN (n7077),
	   .A2 (_net_6284),
	   .A1 (new_n9520_1_) );
   NOR2_X1 g4278 (
	   .ZN (n7072),
	   .A2 (new_n6940_),
	   .A1 (new_n6939_) );
   NAND2_X1 g4277 (
	   .ZN (n7067),
	   .A2 (new_n11006_),
	   .A1 (new_n11001_) );
   AND4_X1 g4276 (
	   .ZN (new_n11006_),
	   .A4 (new_n11005_),
	   .A3 (new_n11004_),
	   .A2 (new_n11003_),
	   .A1 (new_n11002_) );
   NAND2_X1 g4275 (
	   .ZN (new_n11005_),
	   .A2 (_net_6122),
	   .A1 (new_n7209_) );
   NAND2_X1 g4274 (
	   .ZN (new_n11004_),
	   .A2 (new_n7202_),
	   .A1 (new_n9025_1_) );
   NAND2_X1 g4273 (
	   .ZN (new_n11003_),
	   .A2 (new_n7587_),
	   .A1 (new_n7579_) );
   NAND2_X1 g4272 (
	   .ZN (new_n11002_),
	   .A2 (new_n7585_),
	   .A1 (new_n7565_) );
   AND4_X1 g4271 (
	   .ZN (new_n11001_),
	   .A4 (new_n11000_),
	   .A3 (new_n10999_),
	   .A2 (new_n10998_),
	   .A1 (new_n10997_) );
   NAND4_X1 g4270 (
	   .ZN (new_n11000_),
	   .A4 (new_n7194_1_),
	   .A3 (net_6756),
	   .A2 (_net_6822),
	   .A1 (new_n7559_) );
   NAND4_X1 g4269 (
	   .ZN (new_n10999_),
	   .A4 (new_n7191_),
	   .A3 (_net_6822),
	   .A2 (net_6788),
	   .A1 (new_n7560_) );
   NAND3_X1 g4268 (
	   .ZN (new_n10998_),
	   .A3 (new_n7189_),
	   .A2 (net_6820),
	   .A1 (new_n7555_) );
   NAND3_X1 g4267 (
	   .ZN (new_n10997_),
	   .A3 (new_n7196_),
	   .A2 (net_6724),
	   .A1 (new_n7556_) );
   CLKBUF_X1 g4266 (
	   .Z (n7062),
	   .A (_net_7804) );
   OAI21_X1 g4265 (
	   .ZN (n7058),
	   .B2 (new_n6957_1_),
	   .B1 (new_n10994_),
	   .A (new_n10993_) );
   INV_X1 g4264 (
	   .ZN (new_n10994_),
	   .A (_net_7268) );
   NAND2_X1 g4263 (
	   .ZN (new_n10993_),
	   .A2 (new_n7335_1_),
	   .A1 (new_n6949_) );
   MUX2_X1 g4262 (
	   .Z (n7053),
	   .S (new_n10364_),
	   .B (_net_7579),
	   .A (n1163) );
   CLKBUF_X1 g4261 (
	   .Z (n7049),
	   .A (net_6393) );
   CLKBUF_X1 g4260 (
	   .Z (n7045),
	   .A (_net_6182) );
   CLKBUF_X1 g4259 (
	   .Z (n7041),
	   .A (net_6889) );
   CLKBUF_X1 g4258 (
	   .Z (n7036),
	   .A (net_6388) );
   OAI21_X1 g4257 (
	   .ZN (n7032),
	   .B2 (new_n7258_),
	   .B1 (new_n10986_),
	   .A (new_n10985_) );
   INV_X1 g4256 (
	   .ZN (new_n10986_),
	   .A (_net_7298) );
   NAND2_X1 g4255 (
	   .ZN (new_n10985_),
	   .A2 (new_n7321_1_),
	   .A1 (new_n7251_) );
   CLKBUF_X1 g4254 (
	   .Z (n7027),
	   .A (net_7802) );
   NAND2_X1 g4253 (
	   .ZN (n7023),
	   .A2 (new_n10982_),
	   .A1 (new_n10981_) );
   AOI22_X1 g4252 (
	   .ZN (new_n10982_),
	   .B2 (net_7526),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7494) );
   AOI22_X1 g4251 (
	   .ZN (new_n10981_),
	   .B2 (_net_7430),
	   .B1 (new_n7298_),
	   .A2 (net_7462),
	   .A1 (new_n7296_) );
   NAND3_X1 g4250 (
	   .ZN (n7018),
	   .A3 (new_n10979_),
	   .A2 (new_n10978_),
	   .A1 (new_n10974_) );
   AOI22_X1 g4249 (
	   .ZN (new_n10979_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6953),
	   .A2 (new_n10299_),
	   .A1 (new_n6879_) );
   AND3_X1 g4248 (
	   .ZN (new_n10978_),
	   .A3 (new_n10977_),
	   .A2 (new_n10976_),
	   .A1 (new_n10975_) );
   NAND2_X1 g4247 (
	   .ZN (new_n10977_),
	   .A2 (_net_6140),
	   .A1 (new_n6868_) );
   NAND2_X1 g4246 (
	   .ZN (new_n10976_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n9192_1_) );
   NAND2_X1 g4245 (
	   .ZN (new_n10975_),
	   .A2 (new_n6854_),
	   .A1 (new_n9178_1_) );
   AND3_X1 g4244 (
	   .ZN (new_n10974_),
	   .A3 (new_n10973_),
	   .A2 (new_n10972_),
	   .A1 (new_n10971_) );
   NAND4_X1 g4243 (
	   .ZN (new_n10973_),
	   .A4 (new_n6841_),
	   .A3 (net_6921),
	   .A2 (_net_6957),
	   .A1 (new_n6829_) );
   NAND4_X1 g4242 (
	   .ZN (new_n10972_),
	   .A4 (new_n6836_1_),
	   .A3 (_net_6957),
	   .A2 (net_6857),
	   .A1 (new_n6838_) );
   NAND4_X1 g4241 (
	   .ZN (new_n10971_),
	   .A4 (new_n6833_),
	   .A3 (_net_6957),
	   .A2 (net_6889),
	   .A1 (new_n6830_) );
   OAI21_X1 g4240 (
	   .ZN (n7013),
	   .B2 (new_n7652_),
	   .B1 (new_n10969_),
	   .A (new_n10968_) );
   INV_X1 g4239 (
	   .ZN (new_n10969_),
	   .A (_net_7408) );
   NAND2_X1 g4238 (
	   .ZN (new_n10968_),
	   .A2 (new_n8229_),
	   .A1 (new_n7645_) );
   CLKBUF_X1 g4237 (
	   .Z (n7009),
	   .A (net_6597) );
   CLKBUF_X1 g4236 (
	   .Z (n7005),
	   .A (net_6621) );
   MUX2_X1 g4235 (
	   .Z (n7000),
	   .S (new_n7537_),
	   .B (_net_281),
	   .A (_net_7804) );
   OAI21_X1 g4234 (
	   .ZN (n6995),
	   .B2 (new_n6957_1_),
	   .B1 (new_n10963_),
	   .A (new_n10962_) );
   INV_X1 g4233 (
	   .ZN (new_n10963_),
	   .A (_net_7256) );
   NAND2_X1 g4232 (
	   .ZN (new_n10962_),
	   .A2 (new_n8292_),
	   .A1 (new_n6949_) );
   CLKBUF_X1 g4231 (
	   .Z (n6990),
	   .A (_net_7800) );
   CLKBUF_X1 g4230 (
	   .Z (n6986),
	   .A (net_7802) );
   CLKBUF_X1 g4229 (
	   .Z (n6982),
	   .A (_net_6146) );
   CLKBUF_X1 g4228 (
	   .Z (n6977),
	   .A (_net_7816) );
   CLKBUF_X1 g4227 (
	   .Z (n6974),
	   .A (net_7245) );
   OAI221_X1 g4226 (
	   .ZN (n6969),
	   .C2 (new_n7303_),
	   .C1 (new_n10955_),
	   .B2 (new_n7305_),
	   .B1 (new_n7993_),
	   .A (new_n10954_) );
   INV_X1 g4225 (
	   .ZN (new_n10955_),
	   .A (_net_7466) );
   AOI22_X1 g4224 (
	   .ZN (new_n10954_),
	   .B2 (_net_7402),
	   .B1 (new_n9203_),
	   .A2 (_net_7434),
	   .A1 (new_n8694_1_) );
   NAND3_X1 g4223 (
	   .ZN (n6964),
	   .A3 (new_n10952_),
	   .A2 (new_n10951_),
	   .A1 (new_n10947_) );
   AOI22_X1 g4222 (
	   .ZN (new_n10952_),
	   .B2 (new_n7136_),
	   .B1 (net_6681),
	   .A2 (new_n10181_),
	   .A1 (new_n7013_1_) );
   AND3_X1 g4221 (
	   .ZN (new_n10951_),
	   .A3 (new_n10950_),
	   .A2 (new_n10949_),
	   .A1 (new_n10948_) );
   NAND2_X1 g4220 (
	   .ZN (new_n10950_),
	   .A2 (_net_6098),
	   .A1 (new_n6984_) );
   NAND2_X1 g4219 (
	   .ZN (new_n10949_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n7134_) );
   NAND2_X1 g4218 (
	   .ZN (new_n10948_),
	   .A2 (new_n6980_),
	   .A1 (new_n7126_) );
   AND3_X1 g4217 (
	   .ZN (new_n10947_),
	   .A3 (new_n10946_),
	   .A2 (new_n10945_),
	   .A1 (new_n10944_) );
   NAND4_X1 g4216 (
	   .ZN (new_n10946_),
	   .A4 (new_n6987_),
	   .A3 (net_6649),
	   .A2 (_net_6687),
	   .A1 (new_n7114_) );
   NAND4_X1 g4215 (
	   .ZN (new_n10945_),
	   .A4 (new_n6990_1_),
	   .A3 (net_6585),
	   .A2 (_net_6687),
	   .A1 (new_n7118_) );
   NAND4_X1 g4214 (
	   .ZN (new_n10944_),
	   .A4 (new_n6989_),
	   .A3 (net_6617),
	   .A2 (_net_6687),
	   .A1 (new_n7115_) );
   CLKBUF_X1 g4213 (
	   .Z (n6960),
	   .A (_net_7812) );
   CLKBUF_X1 g4212 (
	   .Z (n6957),
	   .A (net_6587) );
   OAI21_X1 g4211 (
	   .ZN (n6952),
	   .B2 (new_n7736_),
	   .B1 (new_n10940_),
	   .A (new_n10939_) );
   INV_X1 g4210 (
	   .ZN (new_n10940_),
	   .A (_net_7500) );
   NAND2_X1 g4209 (
	   .ZN (new_n10939_),
	   .A2 (new_n8066_),
	   .A1 (new_n7732_1_) );
   CLKBUF_X1 g4208 (
	   .Z (n6947),
	   .A (net_6390) );
   MUX2_X1 g4207 (
	   .Z (n6943),
	   .S (new_n7029_),
	   .B (_net_7589),
	   .A (new_n7542_) );
   MUX2_X1 g4206 (
	   .Z (n6938),
	   .S (_net_154),
	   .B (net_310),
	   .A (_net_114) );
   CLKBUF_X1 g4205 (
	   .Z (n6934),
	   .A (net_7150) );
   NAND2_X1 g4204 (
	   .ZN (n6929),
	   .A2 (new_n10933_),
	   .A1 (new_n10932_) );
   AOI22_X1 g4203 (
	   .ZN (new_n10933_),
	   .B2 (new_n6751_),
	   .B1 (_net_7566),
	   .A2 (_net_7662),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g4202 (
	   .ZN (new_n10932_),
	   .B2 (_net_7630),
	   .B1 (new_n8009_),
	   .A2 (new_n7350_),
	   .A1 (_net_7598) );
   OAI21_X1 g4201 (
	   .ZN (n6924),
	   .B2 (new_n7279_),
	   .B1 (new_n10930_),
	   .A (new_n10929_) );
   INV_X1 g4200 (
	   .ZN (new_n10930_),
	   .A (_net_7443) );
   NAND2_X1 g4199 (
	   .ZN (new_n10929_),
	   .A2 (new_n9804_),
	   .A1 (new_n7271_) );
   NOR2_X1 g4198 (
	   .ZN (n6919),
	   .A2 (new_n8104_),
	   .A1 (new_n8675_) );
   NAND2_X1 g4197 (
	   .ZN (n6915),
	   .A2 (new_n10926_),
	   .A1 (new_n10925_) );
   AOI22_X1 g4196 (
	   .ZN (new_n10926_),
	   .B2 (net_7519),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7487) );
   AOI22_X1 g4195 (
	   .ZN (new_n10925_),
	   .B2 (_net_7423),
	   .B1 (new_n7298_),
	   .A2 (net_7455),
	   .A1 (new_n7296_) );
   CLKBUF_X1 g4194 (
	   .Z (n6910),
	   .A (_net_7818) );
   CLKBUF_X1 g4193 (
	   .Z (n6906),
	   .A (_net_7804) );
   CLKBUF_X1 g4192 (
	   .Z (n6902),
	   .A (net_6395) );
   CLKBUF_X1 g4191 (
	   .Z (n6899),
	   .A (net_6607) );
   CLKBUF_X1 g4190 (
	   .Z (n6895),
	   .A (net_7009) );
   AOI21_X1 g4189 (
	   .ZN (n6890),
	   .B2 (new_n7739_),
	   .B1 (new_n10918_),
	   .A (new_n10917_) );
   INV_X1 g4188 (
	   .ZN (new_n10918_),
	   .A (_net_7427) );
   NOR2_X1 g4187 (
	   .ZN (new_n10917_),
	   .A2 (n1173),
	   .A1 (new_n7738_) );
   CLKBUF_X1 g4186 (
	   .Z (n6886),
	   .A (net_6712) );
   NAND3_X1 g4185 (
	   .ZN (n6881),
	   .A3 (new_n10914_),
	   .A2 (new_n10913_),
	   .A1 (new_n10909_) );
   AOI22_X1 g4184 (
	   .ZN (new_n10914_),
	   .B2 (new_n8180_),
	   .B1 (net_7089),
	   .A2 (new_n9972_),
	   .A1 (new_n7060_) );
   AND3_X1 g4183 (
	   .ZN (new_n10913_),
	   .A3 (new_n10912_),
	   .A2 (new_n10911_),
	   .A1 (new_n10910_) );
   NAND2_X1 g4182 (
	   .ZN (new_n10912_),
	   .A2 (_net_6161),
	   .A1 (new_n7091_) );
   NAND2_X1 g4181 (
	   .ZN (new_n10911_),
	   .A2 (new_n7070_),
	   .A1 (new_n8535_1_) );
   NAND2_X1 g4180 (
	   .ZN (new_n10910_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n8521_) );
   AND3_X1 g4179 (
	   .ZN (new_n10909_),
	   .A3 (new_n10908_),
	   .A2 (new_n10907_),
	   .A1 (new_n10906_) );
   NAND4_X1 g4178 (
	   .ZN (new_n10908_),
	   .A4 (new_n7044_),
	   .A3 (_net_7092),
	   .A2 (net_7057),
	   .A1 (new_n8154_) );
   NAND4_X1 g4177 (
	   .ZN (new_n10907_),
	   .A4 (new_n7052_),
	   .A3 (net_6993),
	   .A2 (_net_7092),
	   .A1 (new_n8158_) );
   NAND4_X1 g4176 (
	   .ZN (new_n10906_),
	   .A4 (new_n7050_),
	   .A3 (net_7025),
	   .A2 (_net_7092),
	   .A1 (new_n8155_) );
   CLKBUF_X1 g4175 (
	   .Z (n6876),
	   .A (net_7807) );
   NAND2_X1 g4174 (
	   .ZN (n6872),
	   .A2 (new_n10903_),
	   .A1 (new_n10902_) );
   AOI22_X1 g4173 (
	   .ZN (new_n10903_),
	   .B2 (net_7520),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7488) );
   AOI22_X1 g4172 (
	   .ZN (new_n10902_),
	   .B2 (_net_7424),
	   .B1 (new_n7298_),
	   .A2 (net_7456),
	   .A1 (new_n7296_) );
   CLKBUF_X1 g4171 (
	   .Z (n6867),
	   .A (_net_7823) );
   CLKBUF_X1 g4170 (
	   .Z (n6863),
	   .A (_net_7796) );
   CLKBUF_X1 g4169 (
	   .Z (n6860),
	   .A (net_6470) );
   MUX2_X1 g4168 (
	   .Z (n6855),
	   .S (new_n7436_),
	   .B (_net_5990),
	   .A (net_7799) );
   NAND2_X1 g4167 (
	   .ZN (n6850),
	   .A2 (new_n10896_),
	   .A1 (new_n10895_) );
   AOI22_X1 g4166 (
	   .ZN (new_n10896_),
	   .B2 (new_n6751_),
	   .B1 (_net_7562),
	   .A2 (_net_7658),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g4165 (
	   .ZN (new_n10895_),
	   .B2 (_net_7626),
	   .B1 (new_n8009_),
	   .A2 (new_n7350_),
	   .A1 (_net_7594) );
   OAI21_X1 g4164 (
	   .ZN (n6845),
	   .B2 (new_n7225_),
	   .B1 (new_n10893_),
	   .A (new_n10892_) );
   INV_X1 g4163 (
	   .ZN (new_n10893_),
	   .A (_net_7325) );
   NAND2_X1 g4162 (
	   .ZN (new_n10892_),
	   .A2 (new_n8852_),
	   .A1 (new_n7221_1_) );
   NAND2_X1 g4161 (
	   .ZN (n6840),
	   .A2 (new_n10871_),
	   .A1 (new_n10890_) );
   NAND2_X1 g4160 (
	   .ZN (new_n10890_),
	   .A2 (_net_5960),
	   .A1 (new_n6781_) );
   CLKBUF_X1 g4159 (
	   .Z (n6836),
	   .A (net_7025) );
   MUX2_X1 g4158 (
	   .Z (n6831),
	   .S (new_n7029_),
	   .B (_net_7584),
	   .A (new_n8899_1_) );
   CLKBUF_X1 g4157 (
	   .Z (n6826),
	   .A (_net_7809) );
   CLKBUF_X1 g4156 (
	   .Z (n6822),
	   .A (net_6392) );
   MUX2_X1 g4155 (
	   .Z (n6818),
	   .S (new_n7285_),
	   .B (_net_7700),
	   .A (net_7802) );
   CLKBUF_X1 g4154 (
	   .Z (n6813),
	   .A (_net_7798) );
   CLKBUF_X1 g4153 (
	   .Z (n6809),
	   .A (net_7799) );
   CLKBUF_X1 g4152 (
	   .Z (n6806),
	   .A (net_6990) );
   OAI21_X1 g4151 (
	   .ZN (n6801),
	   .B2 (new_n6957_1_),
	   .B1 (new_n10880_),
	   .A (new_n10879_) );
   INV_X1 g4150 (
	   .ZN (new_n10880_),
	   .A (_net_7258) );
   NAND2_X1 g4149 (
	   .ZN (new_n10879_),
	   .A2 (new_n7495_),
	   .A1 (new_n6949_) );
   CLKBUF_X1 g4148 (
	   .Z (n6796),
	   .A (_net_7801) );
   CLKBUF_X1 g4147 (
	   .Z (n6793),
	   .A (net_7394) );
   OAI21_X1 g4146 (
	   .ZN (n6788),
	   .B2 (new_n7279_),
	   .B1 (new_n10875_),
	   .A (new_n10874_) );
   INV_X1 g4145 (
	   .ZN (new_n10875_),
	   .A (_net_7446) );
   NAND2_X1 g4144 (
	   .ZN (new_n10874_),
	   .A2 (new_n9037_1_),
	   .A1 (new_n7271_) );
   CLKBUF_X1 g4143 (
	   .Z (n6783),
	   .A (_net_7824) );
   AOI21_X1 g4142 (
	   .ZN (n6779),
	   .B2 (new_n10871_),
	   .B1 (new_n10588_),
	   .A (new_n7427_1_) );
   INV_X1 g4141 (
	   .ZN (new_n10871_),
	   .A (_net_5993) );
   NAND2_X1 g4140 (
	   .ZN (n6774),
	   .A2 (new_n10869_),
	   .A1 (new_n10864_) );
   AND4_X1 g4139 (
	   .ZN (new_n10869_),
	   .A4 (new_n10868_),
	   .A3 (new_n10867_),
	   .A2 (new_n10866_),
	   .A1 (new_n10865_) );
   NAND2_X1 g4138 (
	   .ZN (new_n10868_),
	   .A2 (_net_6117),
	   .A1 (new_n7209_) );
   NAND2_X1 g4137 (
	   .ZN (new_n10867_),
	   .A2 (new_n7586_1_),
	   .A1 (new_n10741_) );
   NAND2_X1 g4136 (
	   .ZN (new_n10866_),
	   .A2 (new_n7202_),
	   .A1 (new_n8732_) );
   NAND2_X1 g4135 (
	   .ZN (new_n10865_),
	   .A2 (new_n10830_),
	   .A1 (new_n7565_) );
   AND4_X1 g4134 (
	   .ZN (new_n10864_),
	   .A4 (new_n10863_),
	   .A3 (new_n10862_),
	   .A2 (new_n10861_),
	   .A1 (new_n10860_) );
   NAND4_X1 g4133 (
	   .ZN (new_n10863_),
	   .A4 (new_n7194_1_),
	   .A3 (net_6751),
	   .A2 (_net_6822),
	   .A1 (new_n7559_) );
   NAND4_X1 g4132 (
	   .ZN (new_n10862_),
	   .A4 (new_n7191_),
	   .A3 (_net_6822),
	   .A2 (net_6783),
	   .A1 (new_n7560_) );
   NAND3_X1 g4131 (
	   .ZN (new_n10861_),
	   .A3 (new_n7189_),
	   .A2 (net_6815),
	   .A1 (new_n7555_) );
   NAND3_X1 g4130 (
	   .ZN (new_n10860_),
	   .A3 (new_n7196_),
	   .A2 (net_6719),
	   .A1 (new_n7556_) );
   CLKBUF_X1 g4129 (
	   .Z (n6770),
	   .A (net_6830) );
   NAND3_X1 g4128 (
	   .ZN (n6765),
	   .A3 (new_n10857_),
	   .A2 (new_n10856_),
	   .A1 (new_n10852_) );
   AOI22_X1 g4127 (
	   .ZN (new_n10857_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6949),
	   .A2 (new_n8494_1_),
	   .A1 (new_n6879_) );
   AND3_X1 g4126 (
	   .ZN (new_n10856_),
	   .A3 (new_n10855_),
	   .A2 (new_n10854_),
	   .A1 (new_n10853_) );
   NAND2_X1 g4125 (
	   .ZN (new_n10855_),
	   .A2 (_net_6136),
	   .A1 (new_n6868_) );
   NAND2_X1 g4124 (
	   .ZN (new_n10854_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n8488_) );
   NAND2_X1 g4123 (
	   .ZN (new_n10853_),
	   .A2 (new_n6854_),
	   .A1 (new_n10299_) );
   AND3_X1 g4122 (
	   .ZN (new_n10852_),
	   .A3 (new_n10851_),
	   .A2 (new_n10850_),
	   .A1 (new_n10849_) );
   NAND4_X1 g4121 (
	   .ZN (new_n10851_),
	   .A4 (new_n6841_),
	   .A3 (_net_6957),
	   .A2 (net_6917),
	   .A1 (new_n6829_) );
   NAND4_X1 g4120 (
	   .ZN (new_n10850_),
	   .A4 (new_n6836_1_),
	   .A3 (net_6853),
	   .A2 (_net_6957),
	   .A1 (new_n6838_) );
   NAND4_X1 g4119 (
	   .ZN (new_n10849_),
	   .A4 (new_n6833_),
	   .A3 (_net_6957),
	   .A2 (net_6885),
	   .A1 (new_n6830_) );
   CLKBUF_X1 g4118 (
	   .Z (n6761),
	   .A (net_6728) );
   CLKBUF_X1 g4117 (
	   .Z (n6756),
	   .A (net_6389) );
   CLKBUF_X1 g4116 (
	   .Z (n6752),
	   .A (_net_7794) );
   CLKBUF_X1 g4115 (
	   .Z (n6749),
	   .A (_net_7810) );
   CLKBUF_X1 g4114 (
	   .Z (n6746),
	   .A (net_7549) );
   MUX2_X1 g4113 (
	   .Z (n6741),
	   .S (new_n7504_),
	   .B (_net_7620),
	   .A (new_n8475_) );
   CLKBUF_X1 g4112 (
	   .Z (n6736),
	   .A (net_7799) );
   CLKBUF_X1 g4111 (
	   .Z (n6732),
	   .A (_net_7810) );
   NAND2_X1 g4110 (
	   .ZN (n6727),
	   .A2 (new_n10839_),
	   .A1 (new_n10819_) );
   AND4_X1 g4109 (
	   .ZN (new_n10839_),
	   .A4 (new_n10838_),
	   .A3 (new_n10837_),
	   .A2 (new_n10831_),
	   .A1 (new_n10825_) );
   NAND2_X1 g4108 (
	   .ZN (new_n10838_),
	   .A2 (_net_6113),
	   .A1 (new_n7209_) );
   NAND2_X1 g4107 (
	   .ZN (new_n10837_),
	   .A2 (new_n7587_),
	   .A1 (new_n10836_) );
   NAND4_X1 g4106 (
	   .ZN (new_n10836_),
	   .A4 (new_n10835_),
	   .A3 (new_n10834_),
	   .A2 (new_n10833_),
	   .A1 (new_n10832_) );
   NAND3_X1 g4105 (
	   .ZN (new_n10835_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6797) );
   NAND3_X1 g4104 (
	   .ZN (new_n10834_),
	   .A3 (_net_6824),
	   .A2 (net_6765),
	   .A1 (new_n7186_) );
   NAND3_X1 g4103 (
	   .ZN (new_n10833_),
	   .A3 (_net_6823),
	   .A2 (net_6733),
	   .A1 (new_n7187_) );
   NAND2_X1 g4102 (
	   .ZN (new_n10832_),
	   .A2 (net_6701),
	   .A1 (new_n7566_) );
   NAND2_X1 g4101 (
	   .ZN (new_n10831_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n10830_) );
   NAND4_X1 g4100 (
	   .ZN (new_n10830_),
	   .A4 (new_n10829_),
	   .A3 (new_n10828_),
	   .A2 (new_n10827_),
	   .A1 (new_n10826_) );
   NAND3_X1 g4099 (
	   .ZN (new_n10829_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6799) );
   NAND3_X1 g4098 (
	   .ZN (new_n10828_),
	   .A3 (_net_6824),
	   .A2 (net_6767),
	   .A1 (new_n7186_) );
   NAND3_X1 g4097 (
	   .ZN (new_n10827_),
	   .A3 (_net_6823),
	   .A2 (net_6735),
	   .A1 (new_n7568_) );
   NAND2_X1 g4096 (
	   .ZN (new_n10826_),
	   .A2 (net_6703),
	   .A1 (new_n7566_) );
   NAND2_X1 g4095 (
	   .ZN (new_n10825_),
	   .A2 (new_n10824_),
	   .A1 (new_n7565_) );
   NAND4_X1 g4094 (
	   .ZN (new_n10824_),
	   .A4 (new_n10823_),
	   .A3 (new_n10822_),
	   .A2 (new_n10821_),
	   .A1 (new_n10820_) );
   NAND3_X1 g4093 (
	   .ZN (new_n10823_),
	   .A3 (net_6795),
	   .A2 (_net_6824),
	   .A1 (_net_6823) );
   NAND3_X1 g4092 (
	   .ZN (new_n10822_),
	   .A3 (_net_6824),
	   .A2 (net_6763),
	   .A1 (new_n7570_) );
   NAND3_X1 g4091 (
	   .ZN (new_n10821_),
	   .A3 (net_6731),
	   .A2 (_net_6823),
	   .A1 (new_n7568_) );
   NAND2_X1 g4090 (
	   .ZN (new_n10820_),
	   .A2 (net_6699),
	   .A1 (new_n7566_) );
   AND4_X1 g4089 (
	   .ZN (new_n10819_),
	   .A4 (new_n10818_),
	   .A3 (new_n10817_),
	   .A2 (new_n10816_),
	   .A1 (new_n10815_) );
   NAND4_X1 g4088 (
	   .ZN (new_n10818_),
	   .A4 (new_n7194_1_),
	   .A3 (net_6747),
	   .A2 (_net_6822),
	   .A1 (new_n7559_) );
   NAND4_X1 g4087 (
	   .ZN (new_n10817_),
	   .A4 (new_n7191_),
	   .A3 (net_6779),
	   .A2 (_net_6822),
	   .A1 (new_n7560_) );
   NAND3_X1 g4086 (
	   .ZN (new_n10816_),
	   .A3 (new_n7189_),
	   .A2 (net_6811),
	   .A1 (new_n7555_) );
   NAND3_X1 g4085 (
	   .ZN (new_n10815_),
	   .A3 (new_n7196_),
	   .A2 (net_6715),
	   .A1 (new_n7556_) );
   CLKBUF_X1 g4084 (
	   .Z (n6717),
	   .A (_net_7796) );
   CLKBUF_X1 g4083 (
	   .Z (n6713),
	   .A (_net_7793) );
   AOI21_X1 g4082 (
	   .ZN (n6709),
	   .B2 (new_n7326_1_),
	   .B1 (new_n10811_),
	   .A (new_n10810_) );
   INV_X1 g4081 (
	   .ZN (new_n10811_),
	   .A (_net_7279) );
   NOR2_X1 g4080 (
	   .ZN (new_n10810_),
	   .A2 (n1034),
	   .A1 (new_n7325_) );
   CLKBUF_X1 g4079 (
	   .Z (n6704),
	   .A (_net_7794) );
   CLKBUF_X1 g4078 (
	   .Z (n6700),
	   .A (_net_6157) );
   MUX2_X1 g4077 (
	   .Z (n6695),
	   .S (new_n7504_),
	   .B (_net_7623),
	   .A (new_n9509_) );
   NAND3_X1 g4076 (
	   .ZN (n6691),
	   .A3 (new_n10805_),
	   .A2 (new_n10804_),
	   .A1 (new_n10795_) );
   NAND4_X1 g4075 (
	   .ZN (new_n10805_),
	   .A4 (_net_7696),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR3_X1 g4074 (
	   .ZN (new_n10804_),
	   .A3 (new_n10803_),
	   .A2 (new_n10799_),
	   .A1 (new_n10796_) );
   NAND3_X1 g4073 (
	   .ZN (new_n10803_),
	   .A3 (new_n10802_),
	   .A2 (new_n10801_),
	   .A1 (new_n10800_) );
   NAND4_X1 g4072 (
	   .ZN (new_n10802_),
	   .A4 (net_161),
	   .A3 (x1231),
	   .A2 (new_n7394_),
	   .A1 (new_n7392_) );
   NAND3_X1 g4071 (
	   .ZN (new_n10801_),
	   .A3 (net_198),
	   .A2 (new_n7388_),
	   .A1 (new_n7386_1_) );
   NAND3_X1 g4070 (
	   .ZN (new_n10800_),
	   .A3 (net_235),
	   .A2 (new_n7382_),
	   .A1 (new_n7380_) );
   OAI22_X1 g4069 (
	   .ZN (new_n10799_),
	   .B2 (new_n7378_),
	   .B1 (new_n10798_),
	   .A2 (new_n10797_),
	   .A1 (new_n7374_) );
   INV_X1 g4068 (
	   .ZN (new_n10798_),
	   .A (_net_7725) );
   INV_X1 g4067 (
	   .ZN (new_n10797_),
	   .A (_net_119) );
   AND4_X1 g4066 (
	   .ZN (new_n10796_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7369_),
	   .A1 (_net_6033) );
   NOR2_X1 g4065 (
	   .ZN (new_n10795_),
	   .A2 (new_n10794_),
	   .A1 (new_n10793_) );
   NOR2_X1 g4064 (
	   .ZN (new_n10794_),
	   .A2 (new_n7629_),
	   .A1 (new_n7366_) );
   NOR2_X1 g4063 (
	   .ZN (new_n10793_),
	   .A2 (new_n10792_),
	   .A1 (new_n7362_) );
   INV_X1 g4062 (
	   .ZN (new_n10792_),
	   .A (_net_272) );
   CLKBUF_X1 g4061 (
	   .Z (n6687),
	   .A (net_6997) );
   MUX2_X1 g4060 (
	   .Z (n6682),
	   .S (new_n7538_),
	   .B (_net_278),
	   .A (_net_7801) );
   CLKBUF_X1 g4059 (
	   .Z (n6678),
	   .A (net_6708) );
   CLKBUF_X1 g4058 (
	   .Z (n6674),
	   .A (net_6834) );
   CLKBUF_X1 g4057 (
	   .Z (n6669),
	   .A (net_6390) );
   NAND4_X1 g4056 (
	   .ZN (n6665),
	   .A4 (new_n10785_),
	   .A3 (new_n10784_),
	   .A2 (new_n10780_),
	   .A1 (new_n10774_) );
   NAND2_X1 g4055 (
	   .ZN (new_n10785_),
	   .A2 (new_n6879_),
	   .A1 (new_n8298_) );
   NAND2_X1 g4054 (
	   .ZN (new_n10784_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n10783_) );
   NAND2_X1 g4053 (
	   .ZN (new_n10783_),
	   .A2 (new_n10782_),
	   .A1 (new_n10781_) );
   AOI22_X1 g4052 (
	   .ZN (new_n10782_),
	   .B2 (net_6832),
	   .B1 (new_n6836_1_),
	   .A2 (net_6864),
	   .A1 (new_n6833_) );
   AOI22_X1 g4051 (
	   .ZN (new_n10781_),
	   .B2 (net_6928),
	   .B1 (new_n6873_),
	   .A2 (new_n6841_),
	   .A1 (net_6896) );
   NAND2_X1 g4050 (
	   .ZN (new_n10780_),
	   .A2 (new_n10779_),
	   .A1 (new_n9255_) );
   NAND4_X1 g4049 (
	   .ZN (new_n10779_),
	   .A4 (new_n10778_),
	   .A3 (new_n10777_),
	   .A2 (new_n10776_),
	   .A1 (new_n10775_) );
   NAND3_X1 g4048 (
	   .ZN (new_n10778_),
	   .A3 (_net_6958),
	   .A2 (_net_6959),
	   .A1 (net_6942) );
   NAND3_X1 g4047 (
	   .ZN (new_n10777_),
	   .A3 (net_6910),
	   .A2 (_net_6959),
	   .A1 (new_n6848_) );
   NAND3_X1 g4046 (
	   .ZN (new_n10776_),
	   .A3 (_net_6958),
	   .A2 (net_6878),
	   .A1 (new_n6846_) );
   NAND2_X1 g4045 (
	   .ZN (new_n10775_),
	   .A2 (net_6846),
	   .A1 (new_n6844_) );
   AOI22_X1 g4044 (
	   .ZN (new_n10774_),
	   .B2 (new_n6869_),
	   .B1 (_net_6129),
	   .A2 (new_n6854_),
	   .A1 (new_n6876_1_) );
   CLKBUF_X1 g4043 (
	   .Z (n6661),
	   .A (net_6424) );
   AND2_X1 g4042 (
	   .ZN (n6656),
	   .A2 (net_376),
	   .A1 (new_n7747_) );
   MUX2_X1 g4041 (
	   .Z (n6652),
	   .S (_net_154),
	   .B (net_320),
	   .A (_net_124) );
   CLKBUF_X1 g4040 (
	   .Z (n6648),
	   .A (net_7145) );
   CLKBUF_X1 g4039 (
	   .Z (n6638),
	   .A (_net_7817) );
   NAND4_X1 g4038 (
	   .ZN (n6634),
	   .A4 (new_n10767_),
	   .A3 (new_n10766_),
	   .A2 (new_n10765_),
	   .A1 (new_n10764_) );
   AOI22_X1 g4037 (
	   .ZN (new_n10767_),
	   .B2 (_net_6170),
	   .B1 (new_n7694_),
	   .A2 (new_n7690_),
	   .A1 (new_n9787_1_) );
   NAND2_X1 g4036 (
	   .ZN (new_n10766_),
	   .A2 (new_n7701_),
	   .A1 (new_n8022_) );
   NAND2_X1 g4035 (
	   .ZN (new_n10765_),
	   .A2 (new_n7837_),
	   .A1 (new_n8030_) );
   NAND2_X1 g4034 (
	   .ZN (new_n10764_),
	   .A2 (new_n7832_),
	   .A1 (new_n8026_) );
   CLKBUF_X1 g4033 (
	   .Z (n6629),
	   .A (_net_6085) );
   OAI221_X1 g4032 (
	   .ZN (n6624),
	   .C2 (new_n7312_1_),
	   .C1 (new_n8626_),
	   .B2 (new_n7986_),
	   .B1 (new_n8044_),
	   .A (new_n10761_) );
   AOI22_X1 g4031 (
	   .ZN (new_n10761_),
	   .B2 (_net_7262),
	   .B1 (new_n10556_),
	   .A2 (_net_7326),
	   .A1 (new_n10555_) );
   CLKBUF_X1 g4030 (
	   .Z (n6619),
	   .A (_net_7793) );
   CLKBUF_X1 g4029 (
	   .Z (n6615),
	   .A (_net_7817) );
   CLKBUF_X1 g4028 (
	   .Z (n6611),
	   .A (_net_6096) );
   NOR2_X1 g4027 (
	   .ZN (n6606),
	   .A2 (new_n10756_),
	   .A1 (new_n10755_) );
   XNOR2_X1 g4026 (
	   .ZN (new_n10756_),
	   .B (new_n8923_),
	   .A (new_n9537_1_) );
   NAND4_X1 g4025 (
	   .ZN (new_n10755_),
	   .A4 (new_n10754_),
	   .A3 (new_n10753_),
	   .A2 (new_n10752_),
	   .A1 (new_n10751_) );
   NAND3_X1 g4024 (
	   .ZN (new_n10754_),
	   .A3 (new_n7290_),
	   .A2 (new_n10640_),
	   .A1 (new_n7289_) );
   NAND2_X1 g4023 (
	   .ZN (new_n10753_),
	   .A2 (_net_7097),
	   .A1 (new_n7291_) );
   NAND2_X1 g4022 (
	   .ZN (new_n10752_),
	   .A2 (new_n7072_1_),
	   .A1 (new_n8441_) );
   OAI21_X1 g4021 (
	   .ZN (new_n10751_),
	   .B2 (new_n7057_),
	   .B1 (n2270),
	   .A (_net_7092) );
   OAI21_X1 g4020 (
	   .ZN (n6601),
	   .B2 (new_n7279_),
	   .B1 (new_n10749_),
	   .A (new_n10748_) );
   INV_X1 g4019 (
	   .ZN (new_n10749_),
	   .A (_net_7448) );
   NAND2_X1 g4018 (
	   .ZN (new_n10748_),
	   .A2 (new_n7754_),
	   .A1 (new_n7271_) );
   NAND2_X1 g4017 (
	   .ZN (n6596),
	   .A2 (new_n10746_),
	   .A1 (new_n10736_) );
   AND4_X1 g4016 (
	   .ZN (new_n10746_),
	   .A4 (new_n10745_),
	   .A3 (new_n10744_),
	   .A2 (new_n10743_),
	   .A1 (new_n10742_) );
   NAND2_X1 g4015 (
	   .ZN (new_n10745_),
	   .A2 (_net_6119),
	   .A1 (new_n7209_) );
   NAND2_X1 g4014 (
	   .ZN (new_n10744_),
	   .A2 (new_n7587_),
	   .A1 (new_n8732_) );
   NAND2_X1 g4013 (
	   .ZN (new_n10743_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n8744_) );
   NAND2_X1 g4012 (
	   .ZN (new_n10742_),
	   .A2 (new_n10741_),
	   .A1 (new_n7565_) );
   NAND4_X1 g4011 (
	   .ZN (new_n10741_),
	   .A4 (new_n10740_),
	   .A3 (new_n10739_),
	   .A2 (new_n10738_),
	   .A1 (new_n10737_) );
   NAND3_X1 g4010 (
	   .ZN (new_n10740_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6801) );
   NAND3_X1 g4009 (
	   .ZN (new_n10739_),
	   .A3 (_net_6824),
	   .A2 (net_6769),
	   .A1 (new_n7570_) );
   NAND3_X1 g4008 (
	   .ZN (new_n10738_),
	   .A3 (_net_6823),
	   .A2 (net_6737),
	   .A1 (new_n7568_) );
   NAND2_X1 g4007 (
	   .ZN (new_n10737_),
	   .A2 (net_6705),
	   .A1 (new_n7566_) );
   AND4_X1 g4006 (
	   .ZN (new_n10736_),
	   .A4 (new_n10735_),
	   .A3 (new_n10734_),
	   .A2 (new_n10733_),
	   .A1 (new_n10732_) );
   NAND4_X1 g4005 (
	   .ZN (new_n10735_),
	   .A4 (new_n7194_1_),
	   .A3 (net_6753),
	   .A2 (_net_6822),
	   .A1 (new_n7559_) );
   NAND4_X1 g4004 (
	   .ZN (new_n10734_),
	   .A4 (new_n7191_),
	   .A3 (net_6785),
	   .A2 (_net_6822),
	   .A1 (new_n7560_) );
   NAND3_X1 g4003 (
	   .ZN (new_n10733_),
	   .A3 (new_n7189_),
	   .A2 (net_6817),
	   .A1 (new_n7555_) );
   NAND3_X1 g4002 (
	   .ZN (new_n10732_),
	   .A3 (new_n7196_),
	   .A2 (net_6721),
	   .A1 (new_n7556_) );
   OAI221_X1 g4001 (
	   .ZN (n6591),
	   .C2 (new_n7312_1_),
	   .C1 (new_n10730_),
	   .B2 (new_n7986_),
	   .B1 (new_n9594_),
	   .A (new_n10729_) );
   INV_X1 g4000 (
	   .ZN (new_n10730_),
	   .A (_net_7283) );
   AOI22_X1 g3999 (
	   .ZN (new_n10729_),
	   .B2 (_net_7251),
	   .B1 (new_n10556_),
	   .A2 (_net_7315),
	   .A1 (new_n10555_) );
   CLKBUF_X1 g3998 (
	   .Z (n6586),
	   .A (_net_7817) );
   AOI21_X1 g3997 (
	   .ZN (n6583),
	   .B2 (new_n10726_),
	   .B1 (new_n10725_),
	   .A (new_n8265_) );
   NAND3_X1 g3996 (
	   .ZN (new_n10726_),
	   .A3 (_net_6407),
	   .A2 (_net_6405),
	   .A1 (_net_6406) );
   NOR2_X1 g3995 (
	   .ZN (new_n10725_),
	   .A2 (_net_6411),
	   .A1 (new_n8187_) );
   CLKBUF_X1 g3994 (
	   .Z (n6578),
	   .A (net_132) );
   NOR2_X1 g3993 (
	   .ZN (n6574),
	   .A2 (new_n7275_1_),
	   .A1 (new_n8543_) );
   NAND2_X1 g3992 (
	   .ZN (n6570),
	   .A2 (new_n10721_),
	   .A1 (new_n10720_) );
   NAND2_X1 g3991 (
	   .ZN (new_n10721_),
	   .A2 (new_n7070_),
	   .A1 (new_n9746_1_) );
   AOI22_X1 g3990 (
	   .ZN (new_n10720_),
	   .B2 (new_n7092_),
	   .B1 (_net_6146),
	   .A2 (new_n7089_1_),
	   .A1 (new_n7054_) );
   CLKBUF_X1 g3989 (
	   .Z (n6566),
	   .A (net_6381) );
   CLKBUF_X1 g3988 (
	   .Z (n6563),
	   .A (net_6846) );
   MUX2_X1 g3987 (
	   .Z (n6558),
	   .S (new_n7545_),
	   .B (_net_7654),
	   .A (new_n7762_) );
   CLKBUF_X1 g3986 (
	   .Z (n6554),
	   .A (net_6713) );
   CLKBUF_X1 g3985 (
	   .Z (n6550),
	   .A (net_7397) );
   MUX2_X1 g3984 (
	   .Z (n6545),
	   .S (_net_154),
	   .B (net_314),
	   .A (_net_118) );
   NAND2_X1 g3983 (
	   .ZN (n6540),
	   .A2 (new_n10712_),
	   .A1 (new_n10711_) );
   NAND2_X1 g3982 (
	   .ZN (new_n10712_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n9669_) );
   AOI22_X1 g3981 (
	   .ZN (new_n10711_),
	   .B2 (new_n6869_),
	   .B1 (_net_6126),
	   .A2 (new_n6854_),
	   .A1 (new_n9249_) );
   AND2_X1 g3980 (
	   .ZN (n6535),
	   .A2 (net_376),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g3979 (
	   .Z (n6531),
	   .A (net_6385) );
   AOI21_X1 g3978 (
	   .ZN (n6527),
	   .B2 (new_n10707_),
	   .B1 (new_n10706_),
	   .A (x1034) );
   INV_X1 g3977 (
	   .ZN (new_n10707_),
	   .A (_net_5857) );
   NAND3_X1 g3976 (
	   .ZN (new_n10706_),
	   .A3 (net_7773),
	   .A2 (_net_6001),
	   .A1 (n6643) );
   AOI21_X1 g3975 (
	   .ZN (n6643),
	   .B2 (new_n10704_),
	   .B1 (new_n10703_),
	   .A (new_n6983_) );
   AOI21_X1 g3974 (
	   .ZN (new_n10704_),
	   .B2 (new_n10702_),
	   .B1 (new_n10701_),
	   .A (_net_5964) );
   OAI21_X1 g3973 (
	   .ZN (new_n10703_),
	   .B2 (new_n10702_),
	   .B1 (new_n10701_),
	   .A (new_n8419_) );
   INV_X1 g3972 (
	   .ZN (new_n10702_),
	   .A (_net_5966) );
   NOR2_X1 g3971 (
	   .ZN (new_n10701_),
	   .A2 (_net_5999),
	   .A1 (_net_5965) );
   CLKBUF_X1 g3970 (
	   .Z (n6522),
	   .A (x1501) );
   CLKBUF_X1 g3969 (
	   .Z (n6519),
	   .A (net_6866) );
   CLKBUF_X1 g3968 (
	   .Z (n6515),
	   .A (net_6836) );
   CLKBUF_X1 g3967 (
	   .Z (n6511),
	   .A (net_6604) );
   CLKBUF_X1 g3966 (
	   .Z (n6507),
	   .A (net_6563) );
   CLKBUF_X1 g3965 (
	   .Z (n6502),
	   .A (net_7807) );
   CLKBUF_X1 g3964 (
	   .Z (n6498),
	   .A (_net_6159) );
   OAI221_X1 g3963 (
	   .ZN (n6493),
	   .C2 (new_n7306_),
	   .C1 (new_n10692_),
	   .B2 (new_n7303_),
	   .B1 (new_n10691_),
	   .A (new_n10690_) );
   INV_X1 g3962 (
	   .ZN (new_n10692_),
	   .A (_net_7509) );
   INV_X1 g3961 (
	   .ZN (new_n10691_),
	   .A (_net_7477) );
   AOI22_X1 g3960 (
	   .ZN (new_n10690_),
	   .B2 (_net_7413),
	   .B1 (new_n9203_),
	   .A2 (_net_7445),
	   .A1 (new_n8694_1_) );
   CLKBUF_X1 g3959 (
	   .Z (n6489),
	   .A (net_7242) );
   CLKBUF_X1 g3958 (
	   .Z (n6485),
	   .A (net_6462) );
   CLKBUF_X1 g3957 (
	   .Z (n6480),
	   .A (_net_7796) );
   CLKBUF_X1 g3956 (
	   .Z (n6477),
	   .A (net_7148) );
   CLKBUF_X1 g3955 (
	   .Z (n6472),
	   .A (_net_7812) );
   CLKBUF_X1 g3954 (
	   .Z (n6469),
	   .A (net_6980) );
   CLKBUF_X1 g3953 (
	   .Z (n6464),
	   .A (_net_7817) );
   CLKBUF_X1 g3952 (
	   .Z (n6460),
	   .A (_net_6152) );
   OAI21_X1 g3951 (
	   .ZN (n6455),
	   .B2 (new_n6957_1_),
	   .B1 (new_n10680_),
	   .A (new_n10679_) );
   INV_X1 g3950 (
	   .ZN (new_n10680_),
	   .A (_net_7257) );
   NAND2_X1 g3949 (
	   .ZN (new_n10679_),
	   .A2 (new_n9611_1_),
	   .A1 (new_n6949_) );
   NOR3_X1 g3948 (
	   .ZN (n6450),
	   .A3 (new_n10677_),
	   .A2 (new_n6983_),
	   .A1 (new_n10009_) );
   AOI21_X1 g3947 (
	   .ZN (new_n10677_),
	   .B2 (_net_5967),
	   .B1 (net_6691),
	   .A (_net_6692) );
   CLKBUF_X1 g3946 (
	   .Z (n6446),
	   .A (net_6702) );
   CLKBUF_X1 g3945 (
	   .Z (n6441),
	   .A (net_7802) );
   OAI221_X1 g3944 (
	   .ZN (n6432),
	   .C2 (new_n7312_1_),
	   .C1 (new_n10673_),
	   .B2 (new_n7986_),
	   .B1 (new_n9822_),
	   .A (new_n10672_) );
   INV_X1 g3943 (
	   .ZN (new_n10673_),
	   .A (_net_7282) );
   AOI22_X1 g3942 (
	   .ZN (new_n10672_),
	   .B2 (_net_7250),
	   .B1 (new_n10556_),
	   .A2 (_net_7314),
	   .A1 (new_n10555_) );
   NOR2_X1 g3941 (
	   .ZN (n6427),
	   .A2 (new_n8305_),
	   .A1 (new_n7208_) );
   CLKBUF_X1 g3940 (
	   .Z (n6423),
	   .A (net_6382) );
   CLKBUF_X1 g3939 (
	   .Z (n6419),
	   .A (_net_7795) );
   CLKBUF_X1 g3938 (
	   .Z (n6415),
	   .A (_net_7806) );
   OAI21_X1 g3937 (
	   .ZN (n6411),
	   .B2 (new_n7279_),
	   .B1 (new_n10666_),
	   .A (new_n10665_) );
   INV_X1 g3936 (
	   .ZN (new_n10666_),
	   .A (_net_7438) );
   NAND2_X1 g3935 (
	   .ZN (new_n10665_),
	   .A2 (new_n7963_),
	   .A1 (new_n7271_) );
   CLKBUF_X1 g3934 (
	   .Z (n6407),
	   .A (net_6481) );
   CLKBUF_X1 g3933 (
	   .Z (n6403),
	   .A (net_6738) );
   CLKBUF_X1 g3932 (
	   .Z (n6399),
	   .A (net_6398) );
   NAND3_X1 g3931 (
	   .ZN (n6395),
	   .A3 (new_n10660_),
	   .A2 (new_n10659_),
	   .A1 (new_n10650_) );
   AOI22_X1 g3930 (
	   .ZN (new_n10660_),
	   .B2 (new_n7136_),
	   .B1 (net_6684),
	   .A2 (new_n8800_1_),
	   .A1 (new_n7013_1_) );
   AND3_X1 g3929 (
	   .ZN (new_n10659_),
	   .A3 (new_n10658_),
	   .A2 (new_n10657_),
	   .A1 (new_n10656_) );
   NAND2_X1 g3928 (
	   .ZN (new_n10658_),
	   .A2 (_net_6101),
	   .A1 (new_n6984_) );
   NAND2_X1 g3927 (
	   .ZN (new_n10657_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n10547_) );
   NAND2_X1 g3926 (
	   .ZN (new_n10656_),
	   .A2 (new_n6980_),
	   .A1 (new_n10655_) );
   NAND4_X1 g3925 (
	   .ZN (new_n10655_),
	   .A4 (new_n10654_),
	   .A3 (new_n10653_),
	   .A2 (new_n10652_),
	   .A1 (new_n10651_) );
   NAND3_X1 g3924 (
	   .ZN (new_n10654_),
	   .A3 (_net_6689),
	   .A2 (_net_6688),
	   .A1 (net_6672) );
   NAND3_X1 g3923 (
	   .ZN (new_n10653_),
	   .A3 (net_6640),
	   .A2 (_net_6689),
	   .A1 (new_n7004_) );
   NAND3_X1 g3922 (
	   .ZN (new_n10652_),
	   .A3 (_net_6688),
	   .A2 (net_6608),
	   .A1 (new_n7002_) );
   NAND2_X1 g3921 (
	   .ZN (new_n10651_),
	   .A2 (net_6576),
	   .A1 (new_n6973_) );
   AND3_X1 g3920 (
	   .ZN (new_n10650_),
	   .A3 (new_n10649_),
	   .A2 (new_n10648_),
	   .A1 (new_n10647_) );
   NAND4_X1 g3919 (
	   .ZN (new_n10649_),
	   .A4 (new_n6987_),
	   .A3 (_net_6687),
	   .A2 (net_6652),
	   .A1 (new_n7114_) );
   NAND4_X1 g3918 (
	   .ZN (new_n10648_),
	   .A4 (new_n6990_1_),
	   .A3 (_net_6687),
	   .A2 (net_6588),
	   .A1 (new_n7118_) );
   NAND4_X1 g3917 (
	   .ZN (new_n10647_),
	   .A4 (new_n6989_),
	   .A3 (net_6620),
	   .A2 (_net_6687),
	   .A1 (new_n7115_) );
   CLKBUF_X1 g3916 (
	   .Z (n6390),
	   .A (_net_6165) );
   CLKBUF_X1 g3915 (
	   .Z (n6386),
	   .A (net_7117) );
   MUX2_X1 g3914 (
	   .Z (n6381),
	   .S (new_n7545_),
	   .B (_net_7661),
	   .A (new_n7523_) );
   AOI21_X1 g3913 (
	   .ZN (n6371),
	   .B2 (new_n10641_),
	   .B1 (_net_7098),
	   .A (new_n10642_) );
   OAI21_X1 g3912 (
	   .ZN (new_n10642_),
	   .B2 (_net_7098),
	   .B1 (new_n10641_),
	   .A (_net_6028) );
   NOR3_X1 g3911 (
	   .ZN (new_n10641_),
	   .A3 (new_n10640_),
	   .A2 (new_n8700_),
	   .A1 (new_n8439_) );
   INV_X1 g3910 (
	   .ZN (new_n10640_),
	   .A (_net_7097) );
   CLKBUF_X1 g3909 (
	   .Z (n6367),
	   .A (net_6439) );
   OAI21_X1 g3908 (
	   .ZN (n6362),
	   .B2 (new_n7279_),
	   .B1 (new_n10637_),
	   .A (new_n10636_) );
   INV_X1 g3907 (
	   .ZN (new_n10637_),
	   .A (_net_7440) );
   NAND2_X1 g3906 (
	   .ZN (new_n10636_),
	   .A2 (new_n8229_),
	   .A1 (new_n7272_) );
   CLKBUF_X1 g3905 (
	   .Z (n6357),
	   .A (_net_7817) );
   CLKBUF_X1 g3904 (
	   .Z (n6354),
	   .A (net_6747) );
   CLKBUF_X1 g3903 (
	   .Z (n6350),
	   .A (_net_7794) );
   OAI21_X1 g3902 (
	   .ZN (n6346),
	   .B2 (new_n7111_1_),
	   .B1 (new_n8789_),
	   .A (new_n10631_) );
   NAND2_X1 g3901 (
	   .ZN (new_n10631_),
	   .A2 (new_n9611_1_),
	   .A1 (new_n7100_) );
   CLKBUF_X1 g3900 (
	   .Z (n6342),
	   .A (net_6469) );
   NAND3_X1 g3899 (
	   .ZN (n6337),
	   .A3 (new_n10628_),
	   .A2 (new_n10619_),
	   .A1 (new_n10618_) );
   AND3_X1 g3898 (
	   .ZN (new_n10628_),
	   .A3 (new_n10627_),
	   .A2 (new_n10626_),
	   .A1 (new_n10620_) );
   NAND2_X1 g3897 (
	   .ZN (new_n10627_),
	   .A2 (_net_6074),
	   .A1 (new_n6812_) );
   NAND2_X1 g3896 (
	   .ZN (new_n10626_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n10625_) );
   NAND4_X1 g3895 (
	   .ZN (new_n10625_),
	   .A4 (new_n10624_),
	   .A3 (new_n10623_),
	   .A2 (new_n10622_),
	   .A1 (new_n10621_) );
   NAND3_X1 g3894 (
	   .ZN (new_n10624_),
	   .A3 (net_6528),
	   .A2 (_net_6554),
	   .A1 (_net_6553) );
   NAND3_X1 g3893 (
	   .ZN (new_n10623_),
	   .A3 (_net_6554),
	   .A2 (net_6496),
	   .A1 (new_n6789_) );
   NAND3_X1 g3892 (
	   .ZN (new_n10622_),
	   .A3 (net_6464),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   NAND2_X1 g3891 (
	   .ZN (new_n10621_),
	   .A2 (net_6432),
	   .A1 (new_n6785_) );
   NAND2_X1 g3890 (
	   .ZN (new_n10620_),
	   .A2 (new_n7166_),
	   .A1 (new_n9275_) );
   AOI22_X1 g3889 (
	   .ZN (new_n10619_),
	   .B2 (new_n8211_1_),
	   .B1 (new_n6784_),
	   .A2 (new_n6779_1_),
	   .A1 (net_6542) );
   AND3_X1 g3888 (
	   .ZN (new_n10618_),
	   .A3 (new_n10617_),
	   .A2 (new_n10616_),
	   .A1 (new_n10615_) );
   NAND4_X1 g3887 (
	   .ZN (new_n10617_),
	   .A4 (new_n6775_),
	   .A3 (_net_6552),
	   .A2 (net_6510),
	   .A1 (new_n6763_) );
   NAND4_X1 g3886 (
	   .ZN (new_n10616_),
	   .A4 (new_n6770_1_),
	   .A3 (net_6446),
	   .A2 (_net_6552),
	   .A1 (new_n6772_) );
   NAND4_X1 g3885 (
	   .ZN (new_n10615_),
	   .A4 (new_n6767_),
	   .A3 (_net_6552),
	   .A2 (net_6478),
	   .A1 (new_n6764_) );
   CLKBUF_X1 g3884 (
	   .Z (n6332),
	   .A (net_6396) );
   CLKBUF_X1 g3883 (
	   .Z (n6329),
	   .A (net_7161) );
   MUX2_X1 g3882 (
	   .Z (n6324),
	   .S (new_n7436_),
	   .B (_net_6001),
	   .A (net_7807) );
   CLKBUF_X1 g3881 (
	   .Z (n6319),
	   .A (net_389) );
   CLKBUF_X1 g3880 (
	   .Z (n6316),
	   .A (net_7770) );
   OAI21_X1 g3879 (
	   .ZN (n6311),
	   .B2 (new_n10608_),
	   .B1 (new_n10607_),
	   .A (new_n8416_) );
   NAND2_X1 g3878 (
	   .ZN (new_n10608_),
	   .A2 (_net_5963),
	   .A1 (n8472) );
   OAI21_X1 g3877 (
	   .ZN (new_n10607_),
	   .B2 (new_n10606_),
	   .B1 (new_n10605_),
	   .A (new_n9315_) );
   NOR2_X1 g3876 (
	   .ZN (new_n10606_),
	   .A2 (_net_6558),
	   .A1 (new_n7857_) );
   NOR2_X1 g3875 (
	   .ZN (new_n10605_),
	   .A2 (_net_6555),
	   .A1 (new_n7863_1_) );
   CLKBUF_X1 g3874 (
	   .Z (n6306),
	   .A (net_6393) );
   NOR2_X1 g3873 (
	   .ZN (n6302),
	   .A2 (new_n6934_1_),
	   .A1 (new_n8543_) );
   CLKBUF_X1 g3872 (
	   .Z (n6299),
	   .A (net_7130) );
   NOR3_X1 g3871 (
	   .ZN (n6294),
	   .A3 (new_n10600_),
	   .A2 (new_n7449_),
	   .A1 (new_n10599_) );
   NOR2_X1 g3870 (
	   .ZN (new_n10600_),
	   .A2 (_net_7789),
	   .A1 (new_n10598_) );
   AND2_X1 g3869 (
	   .ZN (new_n10599_),
	   .A2 (_net_7789),
	   .A1 (new_n10598_) );
   AND2_X1 g3868 (
	   .ZN (new_n10598_),
	   .A2 (_net_7788),
	   .A1 (new_n10597_) );
   NOR2_X1 g3867 (
	   .ZN (new_n10597_),
	   .A2 (new_n7443_),
	   .A1 (new_n7450_1_) );
   NAND3_X1 g3866 (
	   .ZN (n6290),
	   .A3 (new_n10595_),
	   .A2 (new_n10594_),
	   .A1 (new_n10585_) );
   OR2_X1 g3865 (
	   .ZN (new_n10595_),
	   .A2 (new_n6808_),
	   .A1 (new_n7365_) );
   NOR3_X1 g3864 (
	   .ZN (new_n10594_),
	   .A3 (new_n10593_),
	   .A2 (new_n10589_),
	   .A1 (new_n10586_) );
   NAND3_X1 g3863 (
	   .ZN (new_n10593_),
	   .A3 (new_n10592_),
	   .A2 (new_n10591_),
	   .A1 (new_n10590_) );
   NAND4_X1 g3862 (
	   .ZN (new_n10592_),
	   .A4 (net_159),
	   .A3 (x1231),
	   .A2 (new_n7394_),
	   .A1 (new_n7392_) );
   NAND3_X1 g3861 (
	   .ZN (new_n10591_),
	   .A3 (net_196),
	   .A2 (new_n7388_),
	   .A1 (new_n7386_1_) );
   NAND3_X1 g3860 (
	   .ZN (new_n10590_),
	   .A3 (net_233),
	   .A2 (new_n7382_),
	   .A1 (new_n7380_) );
   OAI22_X1 g3859 (
	   .ZN (new_n10589_),
	   .B2 (new_n7378_),
	   .B1 (new_n10588_),
	   .A2 (new_n10587_),
	   .A1 (new_n7374_) );
   INV_X1 g3858 (
	   .ZN (new_n10588_),
	   .A (_net_7723) );
   INV_X1 g3857 (
	   .ZN (new_n10587_),
	   .A (_net_117) );
   AND4_X1 g3856 (
	   .ZN (new_n10586_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7369_),
	   .A1 (_net_6031) );
   NOR2_X1 g3855 (
	   .ZN (new_n10585_),
	   .A2 (new_n10584_),
	   .A1 (new_n10583_) );
   NOR2_X1 g3854 (
	   .ZN (new_n10584_),
	   .A2 (new_n7106_),
	   .A1 (new_n7362_) );
   NOR2_X1 g3853 (
	   .ZN (new_n10583_),
	   .A2 (new_n10582_),
	   .A1 (new_n9215_1_) );
   INV_X1 g3852 (
	   .ZN (new_n10582_),
	   .A (_net_7694) );
   CLKBUF_X1 g3851 (
	   .Z (n6285),
	   .A (net_146) );
   OAI221_X1 g3850 (
	   .ZN (n6281),
	   .C2 (new_n6920_),
	   .C1 (new_n9581_),
	   .B2 (new_n6917_),
	   .B1 (new_n7337_),
	   .A (new_n10579_) );
   AOI22_X1 g3849 (
	   .ZN (new_n10579_),
	   .B2 (_net_7268),
	   .B1 (new_n10556_),
	   .A2 (_net_7332),
	   .A1 (new_n10555_) );
   CLKBUF_X1 g3848 (
	   .Z (n6276),
	   .A (_net_5964) );
   OAI221_X1 g3847 (
	   .ZN (n6271),
	   .C2 (new_n7312_1_),
	   .C1 (new_n10576_),
	   .B2 (new_n7986_),
	   .B1 (new_n10425_),
	   .A (new_n10575_) );
   INV_X1 g3846 (
	   .ZN (new_n10576_),
	   .A (_net_7293) );
   AOI22_X1 g3845 (
	   .ZN (new_n10575_),
	   .B2 (_net_7261),
	   .B1 (new_n10556_),
	   .A2 (_net_7325),
	   .A1 (new_n10555_) );
   OAI21_X1 g3844 (
	   .ZN (n6266),
	   .B2 (new_n7279_),
	   .B1 (new_n10573_),
	   .A (new_n10572_) );
   INV_X1 g3843 (
	   .ZN (new_n10573_),
	   .A (_net_7434) );
   NAND2_X1 g3842 (
	   .ZN (new_n10572_),
	   .A2 (new_n7991_),
	   .A1 (new_n7272_) );
   CLKBUF_X1 g3841 (
	   .Z (n6261),
	   .A (x1534) );
   CLKBUF_X1 g3840 (
	   .Z (n6258),
	   .A (net_6750) );
   CLKBUF_X1 g3839 (
	   .Z (n6254),
	   .A (net_6697) );
   OAI221_X1 g3838 (
	   .ZN (n6249),
	   .C2 (new_n7303_),
	   .C1 (new_n10567_),
	   .B2 (new_n7305_),
	   .B1 (new_n9694_),
	   .A (new_n10566_) );
   INV_X1 g3837 (
	   .ZN (new_n10567_),
	   .A (_net_7473) );
   AOI22_X1 g3836 (
	   .ZN (new_n10566_),
	   .B2 (_net_7409),
	   .B1 (new_n9203_),
	   .A2 (_net_7441),
	   .A1 (new_n8694_1_) );
   OAI221_X1 g3835 (
	   .ZN (n6244),
	   .C2 (new_n7303_),
	   .C1 (new_n10464_),
	   .B2 (new_n7306_),
	   .B1 (new_n10028_1_),
	   .A (new_n10564_) );
   AOI22_X1 g3834 (
	   .ZN (new_n10564_),
	   .B2 (_net_7418),
	   .B1 (new_n9203_),
	   .A2 (_net_7450),
	   .A1 (new_n8694_1_) );
   CLKBUF_X1 g3833 (
	   .Z (n6239),
	   .A (net_6400) );
   CLKBUF_X1 g3832 (
	   .Z (n6235),
	   .A (net_7799) );
   NAND2_X1 g3831 (
	   .ZN (n6231),
	   .A2 (n4304),
	   .A1 (new_n7422_1_) );
   OAI221_X1 g3830 (
	   .ZN (n6227),
	   .C2 (new_n6920_),
	   .C1 (new_n10559_),
	   .B2 (new_n6917_),
	   .B1 (new_n10558_),
	   .A (new_n10557_) );
   INV_X1 g3829 (
	   .ZN (new_n10559_),
	   .A (net_7376) );
   INV_X1 g3828 (
	   .ZN (new_n10558_),
	   .A (net_7312) );
   AOI22_X1 g3827 (
	   .ZN (new_n10557_),
	   .B2 (_net_7280),
	   .B1 (new_n10556_),
	   .A2 (net_7344),
	   .A1 (new_n10555_) );
   BUF_X4 g3826 (
	   .Z (new_n10556_),
	   .A (new_n6912_) );
   BUF_X4 g3825 (
	   .Z (new_n10555_),
	   .A (new_n6910_1_) );
   NOR2_X1 g3824 (
	   .ZN (n6222),
	   .A2 (new_n7214_),
	   .A1 (new_n7020_) );
   NAND3_X1 g3823 (
	   .ZN (n6218),
	   .A3 (new_n10552_),
	   .A2 (new_n10551_),
	   .A1 (new_n10542_) );
   AOI22_X1 g3822 (
	   .ZN (new_n10552_),
	   .B2 (new_n7136_),
	   .B1 (net_6682),
	   .A2 (new_n7910_),
	   .A1 (new_n7013_1_) );
   AND3_X1 g3821 (
	   .ZN (new_n10551_),
	   .A3 (new_n10550_),
	   .A2 (new_n10549_),
	   .A1 (new_n10548_) );
   NAND2_X1 g3820 (
	   .ZN (new_n10550_),
	   .A2 (_net_6099),
	   .A1 (new_n6985_) );
   NAND2_X1 g3819 (
	   .ZN (new_n10549_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n8800_1_) );
   NAND2_X1 g3818 (
	   .ZN (new_n10548_),
	   .A2 (new_n6980_),
	   .A1 (new_n10547_) );
   NAND4_X1 g3817 (
	   .ZN (new_n10547_),
	   .A4 (new_n10546_),
	   .A3 (new_n10545_),
	   .A2 (new_n10544_),
	   .A1 (new_n10543_) );
   NAND3_X1 g3816 (
	   .ZN (new_n10546_),
	   .A3 (_net_6689),
	   .A2 (net_6670),
	   .A1 (_net_6688) );
   NAND3_X1 g3815 (
	   .ZN (new_n10545_),
	   .A3 (net_6638),
	   .A2 (_net_6689),
	   .A1 (new_n7004_) );
   NAND3_X1 g3814 (
	   .ZN (new_n10544_),
	   .A3 (_net_6688),
	   .A2 (net_6606),
	   .A1 (new_n7002_) );
   NAND2_X1 g3813 (
	   .ZN (new_n10543_),
	   .A2 (net_6574),
	   .A1 (new_n6973_) );
   AND3_X1 g3812 (
	   .ZN (new_n10542_),
	   .A3 (new_n10541_),
	   .A2 (new_n10540_),
	   .A1 (new_n10539_) );
   NAND4_X1 g3811 (
	   .ZN (new_n10541_),
	   .A4 (new_n6987_),
	   .A3 (net_6650),
	   .A2 (_net_6687),
	   .A1 (new_n7118_) );
   NAND4_X1 g3810 (
	   .ZN (new_n10540_),
	   .A4 (new_n6990_1_),
	   .A3 (_net_6687),
	   .A2 (net_6586),
	   .A1 (new_n7118_) );
   NAND4_X1 g3809 (
	   .ZN (new_n10539_),
	   .A4 (new_n6989_),
	   .A3 (net_6618),
	   .A2 (_net_6687),
	   .A1 (new_n7115_) );
   CLKBUF_X1 g3808 (
	   .Z (n6214),
	   .A (net_7385) );
   OAI21_X1 g3807 (
	   .ZN (n6209),
	   .B2 (new_n6957_1_),
	   .B1 (new_n10536_),
	   .A (new_n10535_) );
   INV_X1 g3806 (
	   .ZN (new_n10536_),
	   .A (_net_7254) );
   NAND2_X1 g3805 (
	   .ZN (new_n10535_),
	   .A2 (new_n9002_),
	   .A1 (new_n6949_) );
   CLKBUF_X1 g3804 (
	   .Z (n6204),
	   .A (net_6397) );
   MUX2_X1 g3803 (
	   .Z (n6200),
	   .S (new_n7285_),
	   .B (_net_7693),
	   .A (_net_7795) );
   CLKBUF_X1 g3802 (
	   .Z (n6195),
	   .A (_net_7813) );
   NAND4_X1 g3801 (
	   .ZN (n6191),
	   .A4 (new_n10530_),
	   .A3 (new_n10529_),
	   .A2 (new_n10528_),
	   .A1 (new_n10527_) );
   NAND2_X1 g3800 (
	   .ZN (new_n10530_),
	   .A2 (new_n7060_),
	   .A1 (new_n7417_1_) );
   NAND2_X1 g3799 (
	   .ZN (new_n10529_),
	   .A2 (new_n7070_),
	   .A1 (new_n7413_1_) );
   NAND2_X1 g3798 (
	   .ZN (new_n10528_),
	   .A2 (new_n8521_),
	   .A1 (new_n7073_) );
   AOI22_X1 g3797 (
	   .ZN (new_n10527_),
	   .B2 (new_n7092_),
	   .B1 (_net_6149),
	   .A2 (new_n7089_1_),
	   .A1 (new_n10526_) );
   NAND2_X1 g3796 (
	   .ZN (new_n10526_),
	   .A2 (new_n10525_),
	   .A1 (new_n10524_) );
   AOI22_X1 g3795 (
	   .ZN (new_n10525_),
	   .B2 (net_6969),
	   .B1 (new_n7063_),
	   .A2 (net_7001),
	   .A1 (new_n7049_1_) );
   AOI22_X1 g3794 (
	   .ZN (new_n10524_),
	   .B2 (net_7065),
	   .B1 (new_n7046_),
	   .A2 (new_n7043_),
	   .A1 (net_7033) );
   OAI21_X1 g3793 (
	   .ZN (n6186),
	   .B2 (new_n8301_),
	   .B1 (new_n10522_),
	   .A (new_n10521_) );
   INV_X1 g3792 (
	   .ZN (new_n10522_),
	   .A (_net_6124) );
   NAND2_X1 g3791 (
	   .ZN (new_n10521_),
	   .A2 (new_n6854_),
	   .A1 (new_n9669_) );
   CLKBUF_X1 g3790 (
	   .Z (n6181),
	   .A (_net_6113) );
   CLKBUF_X1 g3789 (
	   .Z (n6176),
	   .A (_net_6105) );
   NAND4_X1 g3788 (
	   .ZN (n6171),
	   .A4 (new_n10517_),
	   .A3 (new_n10516_),
	   .A2 (new_n10515_),
	   .A1 (new_n10514_) );
   AOI22_X1 g3787 (
	   .ZN (new_n10517_),
	   .B2 (_net_6071),
	   .B1 (new_n6813_1_),
	   .A2 (new_n7166_),
	   .A1 (new_n9238_1_) );
   NAND2_X1 g3786 (
	   .ZN (new_n10516_),
	   .A2 (new_n9095_),
	   .A1 (new_n8205_) );
   NAND2_X1 g3785 (
	   .ZN (new_n10515_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n9871_1_) );
   NAND2_X1 g3784 (
	   .ZN (new_n10514_),
	   .A2 (new_n6784_),
	   .A1 (new_n8142_) );
   AND2_X1 g3783 (
	   .ZN (n6166),
	   .A2 (_net_6208),
	   .A1 (new_n9520_1_) );
   CLKBUF_X1 g3782 (
	   .Z (n6161),
	   .A (_net_7816) );
   CLKBUF_X1 g3781 (
	   .Z (n6158),
	   .A (net_6892) );
   AND2_X1 g3780 (
	   .ZN (n6153),
	   .A2 (_net_6292),
	   .A1 (new_n9520_1_) );
   CLKBUF_X1 g3779 (
	   .Z (n6148),
	   .A (_net_7800) );
   CLKBUF_X1 g3778 (
	   .Z (n6145),
	   .A (net_6594) );
   NOR3_X1 g3777 (
	   .ZN (n6140),
	   .A3 (new_n10506_),
	   .A2 (new_n8325_),
	   .A1 (new_n10505_) );
   AOI21_X1 g3776 (
	   .ZN (new_n10506_),
	   .B2 (net_7680),
	   .B1 (_net_264),
	   .A (_net_7681) );
   NOR3_X1 g3775 (
	   .ZN (new_n10505_),
	   .A3 (new_n6741_1_),
	   .A2 (new_n6960_1_),
	   .A1 (new_n6744_) );
   CLKBUF_X1 g3774 (
	   .Z (n6136),
	   .A (net_6384) );
   CLKBUF_X1 g3773 (
	   .Z (n6132),
	   .A (x1479) );
   CLKBUF_X1 g3772 (
	   .Z (n6128),
	   .A (_net_7803) );
   AOI21_X1 g3771 (
	   .ZN (n6124),
	   .B2 (new_n9142_),
	   .B1 (new_n8469_),
	   .A (new_n7428_) );
   NAND3_X1 g3770 (
	   .ZN (n6119),
	   .A3 (new_n10499_),
	   .A2 (new_n10498_),
	   .A1 (new_n10489_) );
   AOI22_X1 g3769 (
	   .ZN (new_n10499_),
	   .B2 (net_7224),
	   .B1 (new_n7844_),
	   .A2 (new_n8362_1_),
	   .A1 (new_n7837_) );
   AND3_X1 g3768 (
	   .ZN (new_n10498_),
	   .A3 (new_n10497_),
	   .A2 (new_n10496_),
	   .A1 (new_n10490_) );
   NAND2_X1 g3767 (
	   .ZN (new_n10497_),
	   .A2 (_net_6181),
	   .A1 (new_n7694_) );
   NAND2_X1 g3766 (
	   .ZN (new_n10496_),
	   .A2 (new_n7701_),
	   .A1 (new_n10495_) );
   NAND4_X1 g3765 (
	   .ZN (new_n10495_),
	   .A4 (new_n10494_),
	   .A3 (new_n10493_),
	   .A2 (new_n10492_),
	   .A1 (new_n10491_) );
   NAND3_X1 g3764 (
	   .ZN (new_n10494_),
	   .A3 (_net_7228),
	   .A2 (net_7210),
	   .A1 (_net_7229) );
   NAND3_X1 g3763 (
	   .ZN (new_n10493_),
	   .A3 (net_7178),
	   .A2 (_net_7229),
	   .A1 (new_n7823_) );
   NAND3_X1 g3762 (
	   .ZN (new_n10492_),
	   .A3 (_net_7228),
	   .A2 (net_7146),
	   .A1 (new_n7821_) );
   NAND2_X1 g3761 (
	   .ZN (new_n10491_),
	   .A2 (net_7114),
	   .A1 (new_n7819_) );
   NAND2_X1 g3760 (
	   .ZN (new_n10490_),
	   .A2 (new_n7690_),
	   .A1 (new_n8553_) );
   AND3_X1 g3759 (
	   .ZN (new_n10489_),
	   .A3 (new_n10488_),
	   .A2 (new_n10487_),
	   .A1 (new_n10486_) );
   NAND4_X1 g3758 (
	   .ZN (new_n10488_),
	   .A4 (new_n7678_),
	   .A3 (net_7192),
	   .A2 (_net_7227),
	   .A1 (new_n7816_) );
   NAND4_X1 g3757 (
	   .ZN (new_n10487_),
	   .A4 (new_n7683_),
	   .A3 (net_7128),
	   .A2 (_net_7227),
	   .A1 (new_n7816_) );
   NAND4_X1 g3756 (
	   .ZN (new_n10486_),
	   .A4 (new_n7681_1_),
	   .A3 (net_7160),
	   .A2 (_net_7227),
	   .A1 (new_n7813_) );
   CLKBUF_X1 g3755 (
	   .Z (n6114),
	   .A (net_7807) );
   AND2_X1 g3754 (
	   .ZN (n6110),
	   .A2 (net_340),
	   .A1 (new_n7102_1_) );
   CLKBUF_X1 g3753 (
	   .Z (n6106),
	   .A (_net_7824) );
   CLKBUF_X1 g3752 (
	   .Z (n6102),
	   .A (_net_7798) );
   CLKBUF_X1 g3751 (
	   .Z (n6098),
	   .A (_net_6139) );
   OAI21_X1 g3750 (
	   .ZN (n6093),
	   .B2 (new_n7652_),
	   .B1 (new_n10479_),
	   .A (new_n10478_) );
   INV_X1 g3749 (
	   .ZN (new_n10479_),
	   .A (_net_7405) );
   NAND2_X1 g3748 (
	   .ZN (new_n10478_),
	   .A2 (new_n8859_),
	   .A1 (new_n7645_) );
   NOR2_X1 g3747 (
	   .ZN (n6088),
	   .A2 (new_n10476_),
	   .A1 (new_n10475_) );
   NAND4_X1 g3746 (
	   .ZN (new_n10476_),
	   .A4 (_net_6409),
	   .A3 (_net_6404),
	   .A2 (new_n9683_1_),
	   .A1 (new_n8185_) );
   NAND4_X1 g3745 (
	   .ZN (new_n10475_),
	   .A4 (_net_6410),
	   .A3 (new_n9304_),
	   .A2 (new_n9682_),
	   .A1 (new_n8183_1_) );
   NAND2_X1 g3744 (
	   .ZN (n6083),
	   .A2 (new_n10473_),
	   .A1 (new_n10472_) );
   AOI22_X1 g3743 (
	   .ZN (new_n10473_),
	   .B2 (_net_7583),
	   .B1 (new_n6755_),
	   .A2 (net_7615),
	   .A1 (new_n6743_) );
   AOI22_X1 g3742 (
	   .ZN (new_n10472_),
	   .B2 (net_7647),
	   .B1 (new_n8009_),
	   .A2 (new_n7970_1_),
	   .A1 (net_7679) );
   CLKBUF_X1 g3741 (
	   .Z (n6078),
	   .A (x1572) );
   AOI21_X1 g3740 (
	   .ZN (n6074),
	   .B2 (new_n10468_),
	   .B1 (_net_6558),
	   .A (new_n10469_) );
   OAI21_X1 g3739 (
	   .ZN (new_n10469_),
	   .B2 (_net_6558),
	   .B1 (new_n10468_),
	   .A (_net_5984) );
   AND3_X1 g3738 (
	   .ZN (new_n10468_),
	   .A3 (_net_6557),
	   .A2 (net_6556),
	   .A1 (_net_5963) );
   CLKBUF_X1 g3737 (
	   .Z (n6069),
	   .A (_net_7800) );
   CLKBUF_X1 g3736 (
	   .Z (n6066),
	   .A (net_6466) );
   OAI21_X1 g3735 (
	   .ZN (n6061),
	   .B2 (new_n6907_),
	   .B1 (new_n10464_),
	   .A (new_n10463_) );
   INV_X1 g3734 (
	   .ZN (new_n10464_),
	   .A (_net_7482) );
   NAND2_X1 g3733 (
	   .ZN (new_n10463_),
	   .A2 (new_n9502_1_),
	   .A1 (new_n6896_) );
   CLKBUF_X1 g3732 (
	   .Z (n6056),
	   .A (_net_7805) );
   NAND3_X1 g3731 (
	   .ZN (n6052),
	   .A3 (new_n10460_),
	   .A2 (new_n10459_),
	   .A1 (new_n10455_) );
   AOI22_X1 g3730 (
	   .ZN (new_n10460_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6945),
	   .A2 (new_n6878_),
	   .A1 (new_n9253_) );
   AND3_X1 g3729 (
	   .ZN (new_n10459_),
	   .A3 (new_n10458_),
	   .A2 (new_n10457_),
	   .A1 (new_n10456_) );
   NAND2_X1 g3728 (
	   .ZN (new_n10458_),
	   .A2 (_net_6132),
	   .A1 (new_n6869_) );
   NAND2_X1 g3727 (
	   .ZN (new_n10457_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n8502_) );
   NAND2_X1 g3726 (
	   .ZN (new_n10456_),
	   .A2 (new_n6854_),
	   .A1 (new_n8494_1_) );
   AND3_X1 g3725 (
	   .ZN (new_n10455_),
	   .A3 (new_n10454_),
	   .A2 (new_n10453_),
	   .A1 (new_n10452_) );
   NAND4_X1 g3724 (
	   .ZN (new_n10454_),
	   .A4 (new_n6841_),
	   .A3 (_net_6957),
	   .A2 (net_6913),
	   .A1 (new_n6838_) );
   NAND4_X1 g3723 (
	   .ZN (new_n10453_),
	   .A4 (new_n6836_1_),
	   .A3 (_net_6957),
	   .A2 (net_6849),
	   .A1 (new_n6838_) );
   NAND4_X1 g3722 (
	   .ZN (new_n10452_),
	   .A4 (new_n6833_),
	   .A3 (_net_6957),
	   .A2 (net_6881),
	   .A1 (new_n6830_) );
   CLKBUF_X1 g3721 (
	   .Z (n6047),
	   .A (_net_6166) );
   CLKBUF_X1 g3720 (
	   .Z (n6043),
	   .A (net_6733) );
   NAND2_X1 g3719 (
	   .ZN (n6038),
	   .A2 (new_n10448_),
	   .A1 (new_n10447_) );
   AOI22_X1 g3718 (
	   .ZN (new_n10448_),
	   .B2 (_net_7573),
	   .B1 (new_n6755_),
	   .A2 (net_7605),
	   .A1 (new_n6743_) );
   AOI22_X1 g3717 (
	   .ZN (new_n10447_),
	   .B2 (net_7637),
	   .B1 (new_n8009_),
	   .A2 (new_n7970_1_),
	   .A1 (net_7669) );
   CLKBUF_X1 g3716 (
	   .Z (n6034),
	   .A (net_7125) );
   NAND3_X1 g3715 (
	   .ZN (n6029),
	   .A3 (new_n10444_),
	   .A2 (new_n10440_),
	   .A1 (new_n10439_) );
   AND3_X1 g3714 (
	   .ZN (new_n10444_),
	   .A3 (new_n10443_),
	   .A2 (new_n10442_),
	   .A1 (new_n10441_) );
   NAND2_X1 g3713 (
	   .ZN (new_n10443_),
	   .A2 (_net_6081),
	   .A1 (new_n6812_) );
   NAND2_X1 g3712 (
	   .ZN (new_n10442_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n7165_) );
   NAND2_X1 g3711 (
	   .ZN (new_n10441_),
	   .A2 (new_n7166_),
	   .A1 (new_n9089_) );
   AOI22_X1 g3710 (
	   .ZN (new_n10440_),
	   .B2 (new_n7172_1_),
	   .B1 (new_n6784_),
	   .A2 (new_n6779_1_),
	   .A1 (net_6549) );
   AND3_X1 g3709 (
	   .ZN (new_n10439_),
	   .A3 (new_n10438_),
	   .A2 (new_n10437_),
	   .A1 (new_n10436_) );
   NAND4_X1 g3708 (
	   .ZN (new_n10438_),
	   .A4 (new_n6775_),
	   .A3 (_net_6552),
	   .A2 (net_6517),
	   .A1 (new_n6763_) );
   NAND4_X1 g3707 (
	   .ZN (new_n10437_),
	   .A4 (new_n6770_1_),
	   .A3 (_net_6552),
	   .A2 (net_6453),
	   .A1 (new_n6772_) );
   NAND4_X1 g3706 (
	   .ZN (new_n10436_),
	   .A4 (new_n6767_),
	   .A3 (_net_6552),
	   .A2 (net_6485),
	   .A1 (new_n6764_) );
   MUX2_X1 g3705 (
	   .Z (n6024),
	   .S (new_n7029_),
	   .B (_net_7596),
	   .A (new_n8151_) );
   CLKBUF_X1 g3704 (
	   .Z (n6019),
	   .A (_net_6118) );
   CLKBUF_X1 g3703 (
	   .Z (n6014),
	   .A (net_5861) );
   CLKBUF_X1 g3702 (
	   .Z (n6009),
	   .A (net_7802) );
   CLKBUF_X1 g3701 (
	   .Z (n6006),
	   .A (net_7115) );
   CLKBUF_X1 g3700 (
	   .Z (n6002),
	   .A (net_7712) );
   NAND2_X1 g3699 (
	   .ZN (n5997),
	   .A2 (new_n10428_),
	   .A1 (new_n10427_) );
   NAND2_X1 g3698 (
	   .ZN (new_n10428_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n9830_) );
   AOI22_X1 g3697 (
	   .ZN (new_n10427_),
	   .B2 (new_n6813_1_),
	   .B1 (_net_6066),
	   .A2 (new_n7166_),
	   .A1 (new_n8199_) );
   OAI21_X1 g3696 (
	   .ZN (n5992),
	   .B2 (new_n7111_1_),
	   .B1 (new_n10425_),
	   .A (new_n10424_) );
   INV_X1 g3695 (
	   .ZN (new_n10425_),
	   .A (_net_7357) );
   NAND2_X1 g3694 (
	   .ZN (new_n10424_),
	   .A2 (new_n8852_),
	   .A1 (new_n7101_) );
   OAI21_X1 g3693 (
	   .ZN (n5987),
	   .B2 (new_n9569_1_),
	   .B1 (new_n10422_),
	   .A (new_n6963_) );
   NOR2_X1 g3692 (
	   .ZN (new_n10422_),
	   .A2 (_net_6410),
	   .A1 (new_n10421_) );
   NOR2_X1 g3691 (
	   .ZN (new_n10421_),
	   .A2 (new_n8267_),
	   .A1 (new_n9306_) );
   OAI221_X1 g3690 (
	   .ZN (n5982),
	   .C2 (new_n10086_),
	   .C1 (new_n7002_),
	   .B2 (new_n10419_),
	   .B1 (new_n6998_),
	   .A (new_n10417_) );
   NAND2_X1 g3689 (
	   .ZN (new_n10419_),
	   .A2 (new_n7135_),
	   .A1 (new_n10418_) );
   OAI21_X1 g3688 (
	   .ZN (new_n10418_),
	   .B2 (new_n6999_),
	   .B1 (new_n7004_),
	   .A (new_n7002_) );
   OAI21_X1 g3687 (
	   .ZN (new_n10417_),
	   .B2 (new_n6987_),
	   .B1 (new_n6989_),
	   .A (new_n8218_) );
   CLKBUF_X1 g3686 (
	   .Z (n5978),
	   .A (net_6618) );
   OAI21_X1 g3685 (
	   .ZN (n5973),
	   .B2 (new_n7111_1_),
	   .B1 (new_n10414_),
	   .A (new_n10413_) );
   INV_X1 g3684 (
	   .ZN (new_n10414_),
	   .A (_net_7360) );
   NAND2_X1 g3683 (
	   .ZN (new_n10413_),
	   .A2 (new_n7531_),
	   .A1 (new_n7101_) );
   CLKBUF_X1 g3682 (
	   .Z (n5968),
	   .A (_net_7821) );
   CLKBUF_X1 g3681 (
	   .Z (n5964),
	   .A (x1557) );
   MUX2_X1 g3680 (
	   .Z (n5960),
	   .S (new_n7436_),
	   .B (_net_6006),
	   .A (_net_7809) );
   CLKBUF_X1 g3679 (
	   .Z (n5955),
	   .A (_net_6079) );
   CLKBUF_X1 g3678 (
	   .Z (n5951),
	   .A (net_6973) );
   CLKBUF_X1 g3677 (
	   .Z (n5947),
	   .A (net_6562) );
   CLKBUF_X1 g3676 (
	   .Z (n5943),
	   .A (net_6887) );
   MUX2_X1 g3675 (
	   .Z (n5938),
	   .S (new_n10364_),
	   .B (_net_7553),
	   .A (new_n8336_) );
   CLKBUF_X1 g3674 (
	   .Z (n5934),
	   .A (net_7127) );
   CLKBUF_X1 g3673 (
	   .Z (n5930),
	   .A (net_6580) );
   MUX2_X1 g3672 (
	   .Z (n5925),
	   .S (new_n6823_),
	   .B (_net_6040),
	   .A (net_7802) );
   CLKBUF_X1 g3671 (
	   .Z (n5920),
	   .A (_net_7795) );
   CLKBUF_X1 g3670 (
	   .Z (n5917),
	   .A (net_6971) );
   CLKBUF_X1 g3669 (
	   .Z (n5912),
	   .A (_net_7811) );
   CLKBUF_X1 g3668 (
	   .Z (n5908),
	   .A (_net_6180) );
   CLKBUF_X1 g3667 (
	   .Z (n5903),
	   .A (net_7790) );
   OAI21_X1 g3666 (
	   .ZN (n5899),
	   .B2 (new_n7652_),
	   .B1 (new_n10395_),
	   .A (new_n10394_) );
   INV_X1 g3665 (
	   .ZN (new_n10395_),
	   .A (_net_7407) );
   NAND2_X1 g3664 (
	   .ZN (new_n10394_),
	   .A2 (new_n7484_),
	   .A1 (new_n7645_) );
   CLKBUF_X1 g3663 (
	   .Z (n5894),
	   .A (net_6391) );
   MUX2_X1 g3662 (
	   .Z (n5890),
	   .S (new_n7538_),
	   .B (_net_283),
	   .A (_net_7806) );
   XNOR2_X1 g3661 (
	   .ZN (n5885),
	   .B (new_n10390_),
	   .A (new_n10389_) );
   NAND2_X1 g3660 (
	   .ZN (new_n10390_),
	   .A2 (net_7231),
	   .A1 (new_n7823_) );
   XNOR2_X1 g3659 (
	   .ZN (new_n10389_),
	   .B (_net_7232),
	   .A (_net_7229) );
   CLKBUF_X1 g3658 (
	   .Z (n5881),
	   .A (net_6720) );
   CLKBUF_X1 g3657 (
	   .Z (n5876),
	   .A (_net_7822) );
   CLKBUF_X1 g3656 (
	   .Z (n5872),
	   .A (_net_6144) );
   AND2_X1 g3655 (
	   .ZN (n5867),
	   .A2 (net_338),
	   .A1 (new_n7102_1_) );
   CLKBUF_X1 g3654 (
	   .Z (n5864),
	   .A (net_7102) );
   CLKBUF_X1 g3653 (
	   .Z (n5860),
	   .A (net_6479) );
   NOR2_X1 g3652 (
	   .ZN (n5855),
	   .A2 (new_n8187_),
	   .A1 (new_n9685_) );
   AOI21_X1 g3651 (
	   .ZN (n5850),
	   .B2 (new_n10380_),
	   .B1 (new_n10379_),
	   .A (new_n7428_) );
   INV_X1 g3650 (
	   .ZN (new_n10380_),
	   .A (net_6036) );
   INV_X1 g3649 (
	   .ZN (new_n10379_),
	   .A (_net_7734) );
   NAND2_X1 g3648 (
	   .ZN (n5845),
	   .A2 (new_n10377_),
	   .A1 (new_n10376_) );
   AOI22_X1 g3647 (
	   .ZN (new_n10377_),
	   .B2 (_net_7581),
	   .B1 (new_n6755_),
	   .A2 (net_7613),
	   .A1 (new_n6743_) );
   AOI22_X1 g3646 (
	   .ZN (new_n10376_),
	   .B2 (net_7645),
	   .B1 (new_n8009_),
	   .A2 (new_n7970_1_),
	   .A1 (net_7677) );
   CLKBUF_X1 g3645 (
	   .Z (n5840),
	   .A (_net_7793) );
   CLKBUF_X1 g3644 (
	   .Z (n5836),
	   .A (net_7802) );
   CLKBUF_X1 g3643 (
	   .Z (n5833),
	   .A (net_6878) );
   OAI221_X1 g3642 (
	   .ZN (n5828),
	   .C2 (new_n7312_1_),
	   .C1 (new_n9458_),
	   .B2 (new_n7986_),
	   .B1 (new_n7497_),
	   .A (new_n10371_) );
   AOI22_X1 g3641 (
	   .ZN (new_n10371_),
	   .B2 (_net_7258),
	   .B1 (new_n6913_),
	   .A2 (_net_7322),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g3640 (
	   .Z (n5824),
	   .A (net_7113) );
   NAND2_X1 g3639 (
	   .ZN (n5819),
	   .A2 (new_n10368_),
	   .A1 (new_n10367_) );
   AOI22_X1 g3638 (
	   .ZN (new_n10368_),
	   .B2 (new_n6751_),
	   .B1 (_net_7569),
	   .A2 (_net_7665),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g3637 (
	   .ZN (new_n10367_),
	   .B2 (_net_7633),
	   .B1 (new_n8009_),
	   .A2 (new_n6743_),
	   .A1 (_net_7601) );
   AND2_X1 g3636 (
	   .ZN (n5814),
	   .A2 (net_382),
	   .A1 (new_n7018_1_) );
   MUX2_X1 g3635 (
	   .Z (n5809),
	   .S (new_n10364_),
	   .B (_net_7561),
	   .A (new_n10112_1_) );
   BUF_X8 g3634 (
	   .Z (new_n10364_),
	   .A (new_n7608_1_) );
   CLKBUF_X1 g3633 (
	   .Z (n5805),
	   .A (net_6437) );
   CLKBUF_X1 g3632 (
	   .Z (n5801),
	   .A (net_7012) );
   CLKBUF_X1 g3631 (
	   .Z (n5796),
	   .A (net_7802) );
   NOR2_X1 g3630 (
	   .ZN (n5792),
	   .A2 (new_n7508_),
	   .A1 (new_n10359_) );
   INV_X1 g3629 (
	   .ZN (new_n10359_),
	   .A (_net_227) );
   CLKBUF_X1 g3628 (
	   .Z (n5787),
	   .A (_net_7814) );
   CLKBUF_X1 g3627 (
	   .Z (n5783),
	   .A (net_6388) );
   CLKBUF_X1 g3626 (
	   .Z (n5779),
	   .A (_net_7812) );
   NAND3_X1 g3625 (
	   .ZN (n5775),
	   .A3 (new_n10354_),
	   .A2 (new_n10353_),
	   .A1 (new_n10349_) );
   AOI22_X1 g3624 (
	   .ZN (new_n10354_),
	   .B2 (new_n8180_),
	   .B1 (net_7082),
	   .A2 (new_n7086_),
	   .A1 (new_n7060_) );
   AND3_X1 g3623 (
	   .ZN (new_n10353_),
	   .A3 (new_n10352_),
	   .A2 (new_n10351_),
	   .A1 (new_n10350_) );
   NAND2_X1 g3622 (
	   .ZN (new_n10352_),
	   .A2 (_net_6154),
	   .A1 (new_n7091_) );
   NAND2_X1 g3621 (
	   .ZN (new_n10351_),
	   .A2 (new_n7070_),
	   .A1 (new_n8845_1_) );
   NAND2_X1 g3620 (
	   .ZN (new_n10350_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n8837_) );
   AND3_X1 g3619 (
	   .ZN (new_n10349_),
	   .A3 (new_n10348_),
	   .A2 (new_n10347_),
	   .A1 (new_n10346_) );
   NAND4_X1 g3618 (
	   .ZN (new_n10348_),
	   .A4 (new_n7044_),
	   .A3 (net_7050),
	   .A2 (_net_7092),
	   .A1 (new_n8154_) );
   NAND4_X1 g3617 (
	   .ZN (new_n10347_),
	   .A4 (new_n7052_),
	   .A3 (_net_7092),
	   .A2 (net_6986),
	   .A1 (new_n8158_) );
   NAND4_X1 g3616 (
	   .ZN (new_n10346_),
	   .A4 (new_n7050_),
	   .A3 (net_7018),
	   .A2 (_net_7092),
	   .A1 (new_n8155_) );
   CLKBUF_X1 g3615 (
	   .Z (n5771),
	   .A (net_6480) );
   CLKBUF_X1 g3614 (
	   .Z (n5767),
	   .A (net_6590) );
   CLKBUF_X1 g3613 (
	   .Z (n5763),
	   .A (net_6560) );
   CLKBUF_X1 g3612 (
	   .Z (n5758),
	   .A (_net_6131) );
   OAI22_X1 g3611 (
	   .ZN (n5753),
	   .B2 (new_n10340_),
	   .B1 (new_n10052_1_),
	   .A2 (new_n10339_),
	   .A1 (new_n10325_) );
   OAI21_X1 g3610 (
	   .ZN (new_n10340_),
	   .B2 (new_n7446_1_),
	   .B1 (new_n7444_),
	   .A (net_6417) );
   XNOR2_X1 g3609 (
	   .ZN (new_n10339_),
	   .B (new_n10052_1_),
	   .A (new_n10051_) );
   OAI21_X1 g3608 (
	   .ZN (n5748),
	   .B2 (new_n10337_),
	   .B1 (new_n10336_),
	   .A (new_n10335_) );
   XNOR2_X1 g3607 (
	   .ZN (new_n10337_),
	   .B (_net_6825),
	   .A (new_n7189_) );
   INV_X1 g3606 (
	   .ZN (new_n10336_),
	   .A (new_n8765_) );
   AOI22_X1 g3605 (
	   .ZN (new_n10335_),
	   .B2 (_net_6825),
	   .B1 (new_n7210_),
	   .A2 (new_n7560_),
	   .A1 (new_n9628_1_) );
   CLKBUF_X1 g3604 (
	   .Z (n5744),
	   .A (net_7244) );
   MUX2_X1 g3603 (
	   .Z (n5739),
	   .S (new_n7436_),
	   .B (_net_5998),
	   .A (_net_7804) );
   CLKBUF_X1 g3602 (
	   .Z (n5735),
	   .A (net_7026) );
   CLKBUF_X1 g3601 (
	   .Z (n5731),
	   .A (net_7107) );
   CLKBUF_X1 g3600 (
	   .Z (n5727),
	   .A (net_6598) );
   MUX2_X1 g3599 (
	   .Z (n5722),
	   .S (new_n7538_),
	   .B (_net_269),
	   .A (_net_7795) );
   CLKBUF_X1 g3598 (
	   .Z (n5717),
	   .A (_net_7796) );
   CLKBUF_X1 g3597 (
	   .Z (n5713),
	   .A (_net_7806) );
   INV_X1 g3596 (
	   .ZN (n5709),
	   .A (new_n10325_) );
   NAND2_X1 g3595 (
	   .ZN (new_n10325_),
	   .A2 (net_6417),
	   .A1 (new_n7447_) );
   CLKBUF_X1 g3594 (
	   .Z (n5704),
	   .A (_net_7810) );
   OAI221_X1 g3593 (
	   .ZN (n5700),
	   .C2 (new_n7312_1_),
	   .C1 (new_n10198_),
	   .B2 (new_n7986_),
	   .B1 (new_n8107_1_),
	   .A (new_n10322_) );
   AOI22_X1 g3592 (
	   .ZN (new_n10322_),
	   .B2 (_net_7263),
	   .B1 (new_n6913_),
	   .A2 (_net_7327),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g3591 (
	   .Z (n5696),
	   .A (net_6609) );
   AND2_X1 g3590 (
	   .ZN (n5691),
	   .A2 (_net_6282),
	   .A1 (new_n9520_1_) );
   CLKBUF_X1 g3589 (
	   .Z (n5686),
	   .A (x1358) );
   CLKBUF_X1 g3588 (
	   .Z (n5682),
	   .A (_net_7795) );
   CLKBUF_X1 g3587 (
	   .Z (n5679),
	   .A (net_6727) );
   MUX2_X1 g3586 (
	   .Z (n5674),
	   .S (new_n7609_),
	   .B (_net_7564),
	   .A (new_n8151_) );
   AOI21_X1 g3585 (
	   .ZN (n5669),
	   .B2 (new_n8191_),
	   .B1 (_net_7380),
	   .A (new_n10314_) );
   OAI21_X1 g3584 (
	   .ZN (new_n10314_),
	   .B2 (_net_7380),
	   .B1 (new_n8191_),
	   .A (_net_267) );
   CLKBUF_X1 g3583 (
	   .Z (n5664),
	   .A (_net_7813) );
   AND3_X1 g3582 (
	   .ZN (n5660),
	   .A3 (new_n7364_),
	   .A2 (_net_7794),
	   .A1 (new_n6822_1_) );
   CLKBUF_X1 g3581 (
	   .Z (n5655),
	   .A (_net_7795) );
   CLKBUF_X1 g3580 (
	   .Z (n5651),
	   .A (_net_7800) );
   CLKBUF_X1 g3579 (
	   .Z (n5648),
	   .A (net_6983) );
   MUX2_X1 g3578 (
	   .Z (n5643),
	   .S (new_n7504_),
	   .B (_net_7634),
	   .A (new_n8001_) );
   AND2_X1 g3577 (
	   .ZN (n5638),
	   .A2 (_net_6204),
	   .A1 (new_n9520_1_) );
   AOI21_X1 g3576 (
	   .ZN (n5633),
	   .B2 (new_n10305_),
	   .B1 (new_n8919_),
	   .A (new_n7428_) );
   INV_X1 g3575 (
	   .ZN (new_n10305_),
	   .A (_net_7736) );
   NAND3_X1 g3574 (
	   .ZN (n5623),
	   .A3 (new_n10303_),
	   .A2 (new_n10302_),
	   .A1 (new_n10293_) );
   AOI22_X1 g3573 (
	   .ZN (new_n10303_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6951),
	   .A2 (new_n8488_),
	   .A1 (new_n6879_) );
   AND3_X1 g3572 (
	   .ZN (new_n10302_),
	   .A3 (new_n10301_),
	   .A2 (new_n10300_),
	   .A1 (new_n10294_) );
   NAND2_X1 g3571 (
	   .ZN (new_n10301_),
	   .A2 (_net_6138),
	   .A1 (new_n6869_) );
   NAND2_X1 g3570 (
	   .ZN (new_n10300_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n10299_) );
   NAND4_X1 g3569 (
	   .ZN (new_n10299_),
	   .A4 (new_n10298_),
	   .A3 (new_n10297_),
	   .A2 (new_n10296_),
	   .A1 (new_n10295_) );
   NAND3_X1 g3568 (
	   .ZN (new_n10298_),
	   .A3 (net_6937),
	   .A2 (_net_6958),
	   .A1 (_net_6959) );
   NAND3_X1 g3567 (
	   .ZN (new_n10297_),
	   .A3 (net_6905),
	   .A2 (_net_6959),
	   .A1 (new_n6848_) );
   NAND3_X1 g3566 (
	   .ZN (new_n10296_),
	   .A3 (_net_6958),
	   .A2 (net_6873),
	   .A1 (new_n6846_) );
   NAND2_X1 g3565 (
	   .ZN (new_n10295_),
	   .A2 (net_6841),
	   .A1 (new_n6844_) );
   NAND2_X1 g3564 (
	   .ZN (new_n10294_),
	   .A2 (new_n6854_),
	   .A1 (new_n9192_1_) );
   AND3_X1 g3563 (
	   .ZN (new_n10293_),
	   .A3 (new_n10292_),
	   .A2 (new_n10291_),
	   .A1 (new_n10290_) );
   NAND4_X1 g3562 (
	   .ZN (new_n10292_),
	   .A4 (new_n6841_),
	   .A3 (net_6919),
	   .A2 (_net_6957),
	   .A1 (new_n6838_) );
   NAND4_X1 g3561 (
	   .ZN (new_n10291_),
	   .A4 (new_n6836_1_),
	   .A3 (_net_6957),
	   .A2 (net_6855),
	   .A1 (new_n6838_) );
   NAND4_X1 g3560 (
	   .ZN (new_n10290_),
	   .A4 (new_n6833_),
	   .A3 (_net_6957),
	   .A2 (net_6887),
	   .A1 (new_n6830_) );
   CLKBUF_X1 g3559 (
	   .Z (n5618),
	   .A (_net_6067) );
   CLKBUF_X1 g3558 (
	   .Z (n5613),
	   .A (_net_7813) );
   CLKBUF_X1 g3557 (
	   .Z (n5610),
	   .A (_net_7796) );
   CLKBUF_X1 g3556 (
	   .Z (n5606),
	   .A (_net_6172) );
   OAI21_X1 g3555 (
	   .ZN (n5601),
	   .B2 (new_n7652_),
	   .B1 (new_n10284_),
	   .A (new_n10283_) );
   INV_X1 g3554 (
	   .ZN (new_n10284_),
	   .A (_net_7420) );
   NAND2_X1 g3553 (
	   .ZN (new_n10283_),
	   .A2 (new_n9901_),
	   .A1 (new_n7646_) );
   NAND3_X1 g3552 (
	   .ZN (n5596),
	   .A3 (new_n10281_),
	   .A2 (new_n10280_),
	   .A1 (new_n10276_) );
   AOI22_X1 g3551 (
	   .ZN (new_n10281_),
	   .B2 (new_n8180_),
	   .B1 (net_7090),
	   .A2 (new_n8662_1_),
	   .A1 (new_n7060_) );
   AND3_X1 g3550 (
	   .ZN (new_n10280_),
	   .A3 (new_n10279_),
	   .A2 (new_n10278_),
	   .A1 (new_n10277_) );
   NAND2_X1 g3549 (
	   .ZN (new_n10279_),
	   .A2 (_net_6162),
	   .A1 (new_n7091_) );
   NAND2_X1 g3548 (
	   .ZN (new_n10278_),
	   .A2 (new_n7088_),
	   .A1 (new_n7080_) );
   NAND2_X1 g3547 (
	   .ZN (new_n10277_),
	   .A2 (new_n7070_),
	   .A1 (new_n8656_) );
   AND3_X1 g3546 (
	   .ZN (new_n10276_),
	   .A3 (new_n10275_),
	   .A2 (new_n10274_),
	   .A1 (new_n10273_) );
   NAND4_X1 g3545 (
	   .ZN (new_n10275_),
	   .A4 (new_n7044_),
	   .A3 (_net_7092),
	   .A2 (net_7058),
	   .A1 (new_n8154_) );
   NAND4_X1 g3544 (
	   .ZN (new_n10274_),
	   .A4 (new_n7052_),
	   .A3 (net_6994),
	   .A2 (_net_7092),
	   .A1 (new_n8158_) );
   NAND4_X1 g3543 (
	   .ZN (new_n10273_),
	   .A4 (new_n7050_),
	   .A3 (net_7026),
	   .A2 (_net_7092),
	   .A1 (new_n8155_) );
   AND2_X1 g3542 (
	   .ZN (n5591),
	   .A2 (net_378),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g3541 (
	   .Z (n5588),
	   .A (net_7235) );
   CLKBUF_X1 g3540 (
	   .Z (n5584),
	   .A (net_7546) );
   MUX2_X1 g3539 (
	   .Z (n5579),
	   .S (new_n7504_),
	   .B (_net_7622),
	   .A (new_n7762_) );
   CLKBUF_X1 g3538 (
	   .Z (n5575),
	   .A (net_6620) );
   OAI21_X1 g3537 (
	   .ZN (n5570),
	   .B2 (new_n7736_),
	   .B1 (new_n10266_),
	   .A (new_n10265_) );
   INV_X1 g3536 (
	   .ZN (new_n10266_),
	   .A (_net_7502) );
   NAND2_X1 g3535 (
	   .ZN (new_n10265_),
	   .A2 (new_n7963_),
	   .A1 (new_n7732_1_) );
   AOI21_X1 g3534 (
	   .ZN (n5565),
	   .B2 (new_n7739_),
	   .B1 (new_n10263_),
	   .A (new_n10262_) );
   INV_X1 g3533 (
	   .ZN (new_n10263_),
	   .A (_net_7430) );
   NOR2_X1 g3532 (
	   .ZN (new_n10262_),
	   .A2 (n6437),
	   .A1 (new_n7738_) );
   AND2_X1 g3531 (
	   .ZN (n6437),
	   .A2 (net_363),
	   .A1 (new_n6898_) );
   CLKBUF_X1 g3530 (
	   .Z (n5560),
	   .A (_net_7824) );
   CLKBUF_X1 g3529 (
	   .Z (n5556),
	   .A (net_6398) );
   NOR2_X1 g3528 (
	   .ZN (n5552),
	   .A2 (new_n9900_),
	   .A1 (new_n7034_) );
   CLKBUF_X1 g3527 (
	   .Z (n5547),
	   .A (_net_7808) );
   MUX2_X1 g3526 (
	   .Z (n5543),
	   .S (new_n7609_),
	   .B (_net_7577),
	   .A (n3015) );
   CLKBUF_X1 g3525 (
	   .Z (n5539),
	   .A (net_6839) );
   AOI21_X1 g3524 (
	   .ZN (n5534),
	   .B2 (new_n10253_),
	   .B1 (new_n10252_),
	   .A (new_n7428_) );
   NAND3_X1 g3523 (
	   .ZN (new_n10253_),
	   .A3 (net_155),
	   .A2 (net_7771),
	   .A1 (new_n8911_) );
   INV_X1 g3522 (
	   .ZN (new_n10252_),
	   .A (_net_7721) );
   AND2_X1 g3521 (
	   .ZN (n5529),
	   .A2 (new_n10250_),
	   .A1 (new_n10249_) );
   INV_X1 g3520 (
	   .ZN (new_n10250_),
	   .A (x837) );
   AOI211_X1 g3519 (
	   .ZN (new_n10249_),
	   .C2 (new_n10248_),
	   .C1 (new_n10247_),
	   .B (new_n8325_),
	   .A (new_n8885_) );
   AOI21_X1 g3518 (
	   .ZN (new_n10248_),
	   .B2 (new_n10246_),
	   .B1 (new_n10245_),
	   .A (_net_263) );
   OAI21_X1 g3517 (
	   .ZN (new_n10247_),
	   .B2 (new_n10246_),
	   .B1 (new_n10245_),
	   .A (new_n10244_) );
   INV_X1 g3516 (
	   .ZN (new_n10246_),
	   .A (_net_266) );
   NOR2_X1 g3515 (
	   .ZN (new_n10245_),
	   .A2 (_net_293),
	   .A1 (_net_265) );
   INV_X1 g3514 (
	   .ZN (new_n10244_),
	   .A (_net_294) );
   OAI211_X1 g3513 (
	   .ZN (n5525),
	   .C2 (new_n7366_),
	   .C1 (new_n10242_),
	   .B (new_n10241_),
	   .A (new_n10240_) );
   INV_X1 g3512 (
	   .ZN (new_n10242_),
	   .A (net_6024) );
   NAND2_X1 g3511 (
	   .ZN (new_n10241_),
	   .A2 (net_153),
	   .A1 (new_n9995_) );
   AOI21_X1 g3510 (
	   .ZN (new_n10240_),
	   .B2 (new_n9729_1_),
	   .B1 (net_261),
	   .A (new_n10239_) );
   OAI22_X1 g3509 (
	   .ZN (new_n10239_),
	   .B2 (new_n10238_),
	   .B1 (new_n7938_),
	   .A2 (new_n10237_),
	   .A1 (new_n7936_) );
   INV_X1 g3508 (
	   .ZN (new_n10238_),
	   .A (net_187) );
   INV_X1 g3507 (
	   .ZN (new_n10237_),
	   .A (net_224) );
   CLKBUF_X1 g3506 (
	   .Z (n5521),
	   .A (net_7018) );
   NAND4_X1 g3505 (
	   .ZN (n5517),
	   .A4 (new_n10234_),
	   .A3 (new_n10233_),
	   .A2 (new_n10232_),
	   .A1 (new_n10231_) );
   NAND4_X1 g3504 (
	   .ZN (new_n10234_),
	   .A4 (net_7709),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   OR2_X1 g3503 (
	   .ZN (new_n10233_),
	   .A2 (new_n7552_),
	   .A1 (new_n7365_) );
   NAND4_X1 g3502 (
	   .ZN (new_n10232_),
	   .A4 (_net_291),
	   .A3 (x1286),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR2_X1 g3501 (
	   .ZN (new_n10231_),
	   .A2 (new_n10230_),
	   .A1 (new_n10229_) );
   AND2_X1 g3500 (
	   .ZN (new_n10230_),
	   .A2 (net_7738),
	   .A1 (new_n7934_) );
   NAND4_X1 g3499 (
	   .ZN (new_n10229_),
	   .A4 (new_n10228_),
	   .A3 (new_n10227_),
	   .A2 (new_n10226_),
	   .A1 (new_n10225_) );
   NAND4_X1 g3498 (
	   .ZN (new_n10228_),
	   .A4 (_net_174),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g3497 (
	   .ZN (new_n10227_),
	   .A3 (_net_211),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g3496 (
	   .ZN (new_n10226_),
	   .A3 (net_248),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   NAND4_X1 g3495 (
	   .ZN (new_n10225_),
	   .A4 (new_n7354_1_),
	   .A3 (net_148),
	   .A2 (x1261),
	   .A1 (new_n7370_) );
   CLKBUF_X1 g3494 (
	   .Z (n5513),
	   .A (net_6024) );
   OAI21_X1 g3493 (
	   .ZN (n5508),
	   .B2 (new_n6907_),
	   .B1 (new_n10222_),
	   .A (new_n10221_) );
   INV_X1 g3492 (
	   .ZN (new_n10222_),
	   .A (_net_7467) );
   NAND2_X1 g3491 (
	   .ZN (new_n10221_),
	   .A2 (new_n9722_),
	   .A1 (new_n6897_) );
   CLKBUF_X1 g3490 (
	   .Z (n5504),
	   .A (net_7100) );
   CLKBUF_X1 g3489 (
	   .Z (n5500),
	   .A (net_6575) );
   MUX2_X1 g3488 (
	   .Z (n5495),
	   .S (new_n7538_),
	   .B (_net_270),
	   .A (_net_7796) );
   OAI21_X1 g3487 (
	   .ZN (n5490),
	   .B2 (new_n7736_),
	   .B1 (new_n10216_),
	   .A (new_n10215_) );
   INV_X1 g3486 (
	   .ZN (new_n10216_),
	   .A (_net_7513) );
   NAND2_X1 g3485 (
	   .ZN (new_n10215_),
	   .A2 (new_n6904_),
	   .A1 (new_n7733_) );
   CLKBUF_X1 g3484 (
	   .Z (n5486),
	   .A (net_387) );
   CLKBUF_X1 g3483 (
	   .Z (n5481),
	   .A (_net_7815) );
   MUX2_X1 g3482 (
	   .Z (n5477),
	   .S (new_n7029_),
	   .B (_net_7587),
	   .A (new_n9197_) );
   AND2_X1 g3481 (
	   .ZN (n5472),
	   .A2 (net_380),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g3480 (
	   .Z (n5469),
	   .A (net_6610) );
   NOR2_X1 g3479 (
	   .ZN (n5464),
	   .A2 (new_n7107_1_),
	   .A1 (new_n8675_) );
   CLKBUF_X1 g3478 (
	   .Z (n5460),
	   .A (_net_6075) );
   MUX2_X1 g3477 (
	   .Z (n5455),
	   .S (new_n7436_),
	   .B (_net_5987),
	   .A (_net_7796) );
   CLKBUF_X1 g3476 (
	   .Z (n5451),
	   .A (net_6436) );
   MUX2_X1 g3475 (
	   .Z (n5446),
	   .S (_net_154),
	   .B (net_315),
	   .A (_net_119) );
   CLKBUF_X1 g3474 (
	   .Z (n5441),
	   .A (_net_7824) );
   CLKBUF_X1 g3473 (
	   .Z (n5437),
	   .A (net_6395) );
   CLKBUF_X1 g3472 (
	   .Z (n5433),
	   .A (_net_7801) );
   MUX2_X1 g3471 (
	   .Z (n5429),
	   .S (new_n6823_),
	   .B (_net_6030),
	   .A (_net_7795) );
   CLKBUF_X1 g3470 (
	   .Z (n5424),
	   .A (_net_7797) );
   OAI21_X1 g3469 (
	   .ZN (n5420),
	   .B2 (new_n7258_),
	   .B1 (new_n10198_),
	   .A (new_n10197_) );
   INV_X1 g3468 (
	   .ZN (new_n10198_),
	   .A (_net_7295) );
   NAND2_X1 g3467 (
	   .ZN (new_n10197_),
	   .A2 (new_n8105_),
	   .A1 (new_n7252_1_) );
   CLKBUF_X1 g3466 (
	   .Z (n5415),
	   .A (_net_7804) );
   MUX2_X1 g3465 (
	   .Z (n5411),
	   .S (new_n7504_),
	   .B (_net_7631),
	   .A (new_n8687_) );
   AOI21_X1 g3464 (
	   .ZN (n5406),
	   .B2 (new_n7739_),
	   .B1 (new_n10193_),
	   .A (new_n10192_) );
   INV_X1 g3463 (
	   .ZN (new_n10193_),
	   .A (_net_7429) );
   NOR2_X1 g3462 (
	   .ZN (new_n10192_),
	   .A2 (n420),
	   .A1 (new_n7738_) );
   CLKBUF_X1 g3461 (
	   .Z (n5402),
	   .A (net_7151) );
   OAI221_X1 g3460 (
	   .ZN (n5397),
	   .C2 (new_n6920_),
	   .C1 (new_n10189_),
	   .B2 (new_n6917_),
	   .B1 (new_n7257_),
	   .A (new_n10188_) );
   INV_X1 g3459 (
	   .ZN (new_n10189_),
	   .A (_net_7349) );
   AOI22_X1 g3458 (
	   .ZN (new_n10188_),
	   .B2 (_net_7253),
	   .B1 (new_n6913_),
	   .A2 (_net_7317),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g3457 (
	   .Z (n5393),
	   .A (net_7021) );
   NAND3_X1 g3456 (
	   .ZN (n5388),
	   .A3 (new_n10185_),
	   .A2 (new_n10184_),
	   .A1 (new_n10175_) );
   AOI22_X1 g3455 (
	   .ZN (new_n10185_),
	   .B2 (new_n7136_),
	   .B1 (net_6679),
	   .A2 (new_n9328_),
	   .A1 (new_n7013_1_) );
   AND3_X1 g3454 (
	   .ZN (new_n10184_),
	   .A3 (new_n10183_),
	   .A2 (new_n10182_),
	   .A1 (new_n10176_) );
   NAND2_X1 g3453 (
	   .ZN (new_n10183_),
	   .A2 (_net_6096),
	   .A1 (new_n6985_) );
   NAND2_X1 g3452 (
	   .ZN (new_n10182_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n10181_) );
   NAND4_X1 g3451 (
	   .ZN (new_n10181_),
	   .A4 (new_n10180_),
	   .A3 (new_n10179_),
	   .A2 (new_n10178_),
	   .A1 (new_n10177_) );
   NAND3_X1 g3450 (
	   .ZN (new_n10180_),
	   .A3 (net_6665),
	   .A2 (_net_6689),
	   .A1 (_net_6688) );
   NAND3_X1 g3449 (
	   .ZN (new_n10179_),
	   .A3 (_net_6689),
	   .A2 (net_6633),
	   .A1 (new_n7004_) );
   NAND3_X1 g3448 (
	   .ZN (new_n10178_),
	   .A3 (net_6601),
	   .A2 (_net_6688),
	   .A1 (new_n7002_) );
   NAND2_X1 g3447 (
	   .ZN (new_n10177_),
	   .A2 (net_6569),
	   .A1 (new_n6973_) );
   NAND2_X1 g3446 (
	   .ZN (new_n10176_),
	   .A2 (new_n6980_),
	   .A1 (new_n7134_) );
   AND3_X1 g3445 (
	   .ZN (new_n10175_),
	   .A3 (new_n10174_),
	   .A2 (new_n10173_),
	   .A1 (new_n10172_) );
   NAND4_X1 g3444 (
	   .ZN (new_n10174_),
	   .A4 (new_n6987_),
	   .A3 (net_6647),
	   .A2 (_net_6687),
	   .A1 (new_n7118_) );
   NAND4_X1 g3443 (
	   .ZN (new_n10173_),
	   .A4 (new_n6990_1_),
	   .A3 (net_6583),
	   .A2 (_net_6687),
	   .A1 (new_n7118_) );
   NAND4_X1 g3442 (
	   .ZN (new_n10172_),
	   .A4 (new_n6989_),
	   .A3 (net_6615),
	   .A2 (_net_6687),
	   .A1 (new_n7115_) );
   CLKBUF_X1 g3441 (
	   .Z (n5383),
	   .A (_net_7819) );
   CLKBUF_X1 g3440 (
	   .Z (n5380),
	   .A (net_6729) );
   CLKBUF_X1 g3439 (
	   .Z (n5375),
	   .A (net_143) );
   MUX2_X1 g3438 (
	   .Z (n5370),
	   .S (new_n7545_),
	   .B (_net_7657),
	   .A (new_n10112_1_) );
   CLKBUF_X1 g3437 (
	   .Z (n5366),
	   .A (net_6860) );
   CLKBUF_X1 g3436 (
	   .Z (n5362),
	   .A (net_6460) );
   CLKBUF_X1 g3435 (
	   .Z (n5358),
	   .A (net_6454) );
   AOI21_X1 g3434 (
	   .ZN (n5353),
	   .B2 (new_n7326_1_),
	   .B1 (new_n10163_),
	   .A (new_n10162_) );
   INV_X1 g3433 (
	   .ZN (new_n10163_),
	   .A (_net_7280) );
   NOR2_X1 g3432 (
	   .ZN (new_n10162_),
	   .A2 (n875),
	   .A1 (new_n7325_) );
   CLKBUF_X1 g3431 (
	   .Z (n5349),
	   .A (net_6987) );
   OAI21_X1 g3430 (
	   .ZN (n5344),
	   .B2 (new_n10159_),
	   .B1 (new_n9434_),
	   .A (new_n10158_1_) );
   NAND2_X1 g3429 (
	   .ZN (new_n10159_),
	   .A2 (new_n9440_),
	   .A1 (n7691) );
   NAND3_X1 g3428 (
	   .ZN (new_n10158_1_),
	   .A3 (new_n10157_),
	   .A2 (new_n9675_),
	   .A1 (new_n9673_1_) );
   OAI21_X1 g3427 (
	   .ZN (new_n10157_),
	   .B2 (new_n9438_),
	   .B1 (new_n9433_),
	   .A (new_n9434_) );
   CLKBUF_X1 g3426 (
	   .Z (n5339),
	   .A (_net_6161) );
   CLKBUF_X1 g3425 (
	   .Z (n5335),
	   .A (net_7002) );
   MUX2_X1 g3424 (
	   .Z (n5330),
	   .S (new_n7545_),
	   .B (_net_7662),
	   .A (new_n9405_1_) );
   CLKBUF_X1 g3423 (
	   .Z (n5326),
	   .A (net_6844) );
   AOI21_X1 g3422 (
	   .ZN (n5321),
	   .B2 (new_n10151_),
	   .B1 (new_n10150_1_),
	   .A (new_n8325_) );
   NAND2_X1 g3421 (
	   .ZN (new_n10151_),
	   .A2 (new_n7502_),
	   .A1 (new_n7026_) );
   OR2_X1 g3420 (
	   .ZN (new_n10150_1_),
	   .A2 (new_n7502_),
	   .A1 (new_n7026_) );
   AOI21_X1 g3419 (
	   .ZN (n5316),
	   .B2 (net_309),
	   .B1 (_net_5985),
	   .A (new_n10148_) );
   NAND3_X1 g3418 (
	   .ZN (new_n10148_),
	   .A3 (_net_5984),
	   .A2 (new_n10147_),
	   .A1 (new_n7655_) );
   INV_X1 g3417 (
	   .ZN (new_n10147_),
	   .A (net_7750) );
   CLKBUF_X1 g3416 (
	   .Z (n5312),
	   .A (net_7006) );
   OAI21_X1 g3415 (
	   .ZN (n5307),
	   .B2 (new_n7652_),
	   .B1 (new_n10144_),
	   .A (new_n10143_) );
   INV_X1 g3414 (
	   .ZN (new_n10144_),
	   .A (_net_7411) );
   NAND2_X1 g3413 (
	   .ZN (new_n10143_),
	   .A2 (new_n9804_),
	   .A1 (new_n7646_) );
   CLKBUF_X1 g3412 (
	   .Z (n5302),
	   .A (_net_6128) );
   CLKBUF_X1 g3411 (
	   .Z (n5298),
	   .A (net_6965) );
   MUX2_X1 g3410 (
	   .Z (n5293),
	   .S (new_n7029_),
	   .B (_net_7599),
	   .A (new_n8687_) );
   CLKBUF_X1 g3409 (
	   .Z (n5288),
	   .A (net_6395) );
   AND2_X1 g3408 (
	   .ZN (n5284),
	   .A2 (_net_6283),
	   .A1 (new_n9520_1_) );
   AOI21_X1 g3407 (
	   .ZN (n5279),
	   .B2 (new_n10136_),
	   .B1 (new_n10135_),
	   .A (new_n7428_) );
   INV_X1 g3406 (
	   .ZN (new_n10136_),
	   .A (_net_7731) );
   INV_X1 g3405 (
	   .ZN (new_n10135_),
	   .A (net_6025) );
   OAI21_X1 g3404 (
	   .ZN (n5274),
	   .B2 (new_n7258_),
	   .B1 (new_n10133_),
	   .A (new_n10132_1_) );
   INV_X1 g3403 (
	   .ZN (new_n10133_),
	   .A (_net_7292) );
   NAND2_X1 g3402 (
	   .ZN (new_n10132_1_),
	   .A2 (new_n10131_),
	   .A1 (new_n7252_1_) );
   OAI21_X1 g3401 (
	   .ZN (new_n10131_),
	   .B2 (new_n10130_),
	   .B1 (new_n6951_),
	   .A (new_n10129_) );
   INV_X1 g3400 (
	   .ZN (new_n10130_),
	   .A (net_7244) );
   AOI22_X1 g3399 (
	   .ZN (new_n10129_),
	   .B2 (net_338),
	   .B1 (_net_269),
	   .A2 (_net_270),
	   .A1 (net_336) );
   CLKBUF_X1 g3398 (
	   .Z (n5269),
	   .A (_net_7798) );
   OAI21_X1 g3397 (
	   .ZN (n5265),
	   .B2 (new_n7652_),
	   .B1 (new_n10126_),
	   .A (new_n10125_) );
   INV_X1 g3396 (
	   .ZN (new_n10126_),
	   .A (_net_7416) );
   NAND2_X1 g3395 (
	   .ZN (new_n10125_),
	   .A2 (new_n7754_),
	   .A1 (new_n7646_) );
   CLKBUF_X1 g3394 (
	   .Z (n5261),
	   .A (net_6843) );
   MUX2_X1 g3393 (
	   .Z (n5256),
	   .S (new_n7609_),
	   .B (_net_7567),
	   .A (new_n8687_) );
   OAI21_X1 g3392 (
	   .ZN (n5251),
	   .B2 (new_n7258_),
	   .B1 (new_n7466_),
	   .A (new_n10121_) );
   NAND2_X1 g3391 (
	   .ZN (new_n10121_),
	   .A2 (new_n9560_),
	   .A1 (new_n7252_1_) );
   CLKBUF_X1 g3390 (
	   .Z (n5246),
	   .A (_net_7797) );
   CLKBUF_X1 g3389 (
	   .Z (n5242),
	   .A (_net_7814) );
   CLKBUF_X1 g3388 (
	   .Z (n5239),
	   .A (net_6487) );
   CLKBUF_X1 g3387 (
	   .Z (n5234),
	   .A (_net_7806) );
   AOI21_X1 g3386 (
	   .ZN (n5230),
	   .B2 (new_n7739_),
	   .B1 (new_n10115_),
	   .A (new_n10114_) );
   INV_X1 g3385 (
	   .ZN (new_n10115_),
	   .A (_net_7422) );
   NOR2_X1 g3384 (
	   .ZN (new_n10114_),
	   .A2 (n5027),
	   .A1 (new_n7738_) );
   MUX2_X1 g3383 (
	   .Z (n5225),
	   .S (new_n7029_),
	   .B (_net_7593),
	   .A (new_n10112_1_) );
   OAI21_X1 g3382 (
	   .ZN (new_n10112_1_),
	   .B2 (new_n10111_),
	   .B1 (new_n7019_),
	   .A (new_n10110_) );
   INV_X1 g3381 (
	   .ZN (new_n10111_),
	   .A (net_7545) );
   AOI22_X1 g3380 (
	   .ZN (new_n10110_),
	   .B2 (_net_292),
	   .B1 (net_375),
	   .A2 (_net_291),
	   .A1 (net_377) );
   CLKBUF_X1 g3379 (
	   .Z (n5221),
	   .A (net_6857) );
   CLKBUF_X1 g3378 (
	   .Z (n5217),
	   .A (net_6569) );
   NAND2_X1 g3377 (
	   .ZN (n5212),
	   .A2 (new_n10106_),
	   .A1 (new_n10101_) );
   AND4_X1 g3376 (
	   .ZN (new_n10106_),
	   .A4 (new_n10105_),
	   .A3 (new_n10104_),
	   .A2 (new_n10103_1_),
	   .A1 (new_n10102_) );
   NAND2_X1 g3375 (
	   .ZN (new_n10105_),
	   .A2 (_net_6114),
	   .A1 (new_n7210_) );
   NAND2_X1 g3374 (
	   .ZN (new_n10104_),
	   .A2 (new_n7587_),
	   .A1 (new_n9493_) );
   NAND2_X1 g3373 (
	   .ZN (new_n10103_1_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n8617_) );
   NAND2_X1 g3372 (
	   .ZN (new_n10102_),
	   .A2 (new_n9032_),
	   .A1 (new_n7565_) );
   AND4_X1 g3371 (
	   .ZN (new_n10101_),
	   .A4 (new_n10100_),
	   .A3 (new_n10099_1_),
	   .A2 (new_n10098_),
	   .A1 (new_n10097_) );
   NAND4_X1 g3370 (
	   .ZN (new_n10100_),
	   .A4 (new_n7194_1_),
	   .A3 (net_6748),
	   .A2 (_net_6822),
	   .A1 (new_n7559_) );
   NAND4_X1 g3369 (
	   .ZN (new_n10099_1_),
	   .A4 (new_n7191_),
	   .A3 (net_6780),
	   .A2 (_net_6822),
	   .A1 (new_n7560_) );
   NAND3_X1 g3368 (
	   .ZN (new_n10098_),
	   .A3 (new_n7189_),
	   .A2 (net_6812),
	   .A1 (new_n7555_) );
   NAND3_X1 g3367 (
	   .ZN (new_n10097_),
	   .A3 (new_n7196_),
	   .A2 (net_6716),
	   .A1 (new_n7556_) );
   OAI221_X1 g3366 (
	   .ZN (n5207),
	   .C2 (new_n10095_),
	   .C1 (new_n8327_),
	   .B2 (new_n10093_),
	   .B1 (new_n10090_),
	   .A (new_n10092_) );
   XNOR2_X1 g3365 (
	   .ZN (new_n10095_),
	   .B (new_n10090_),
	   .A (new_n10094_1_) );
   NAND3_X1 g3364 (
	   .ZN (new_n10094_1_),
	   .A3 (_net_7685),
	   .A2 (_net_7684),
	   .A1 (_net_7683) );
   NAND2_X1 g3363 (
	   .ZN (new_n10093_),
	   .A2 (_net_289),
	   .A1 (new_n7024_) );
   NAND4_X1 g3362 (
	   .ZN (new_n10092_),
	   .A4 (new_n10091_),
	   .A3 (new_n7020_),
	   .A2 (new_n10089_1_),
	   .A1 (new_n8326_) );
   OAI21_X1 g3361 (
	   .ZN (new_n10091_),
	   .B2 (new_n7027_1_),
	   .B1 (new_n7502_),
	   .A (new_n10090_) );
   INV_X1 g3360 (
	   .ZN (new_n10090_),
	   .A (_net_7686) );
   NAND2_X1 g3359 (
	   .ZN (new_n10089_1_),
	   .A2 (_net_7686),
	   .A1 (new_n7543_1_) );
   CLKBUF_X1 g3358 (
	   .Z (n5202),
	   .A (_net_7811) );
   OAI21_X1 g3357 (
	   .ZN (n5198),
	   .B2 (new_n10086_),
	   .B1 (new_n10085_),
	   .A (new_n10084_1_) );
   INV_X1 g3356 (
	   .ZN (new_n10086_),
	   .A (new_n6985_) );
   INV_X1 g3355 (
	   .ZN (new_n10085_),
	   .A (_net_6084) );
   NAND2_X1 g3354 (
	   .ZN (new_n10084_1_),
	   .A2 (new_n6980_),
	   .A1 (new_n7011_) );
   CLKBUF_X1 g3353 (
	   .Z (n5193),
	   .A (net_7802) );
   CLKBUF_X1 g3352 (
	   .Z (n5189),
	   .A (_net_7794) );
   CLKBUF_X1 g3351 (
	   .Z (n5186),
	   .A (net_7691) );
   CLKBUF_X1 g3350 (
	   .Z (n5181),
	   .A (x1519) );
   CLKBUF_X1 g3349 (
	   .Z (n5178),
	   .A (net_6841) );
   CLKBUF_X1 g3348 (
	   .Z (n5173),
	   .A (_net_7808) );
   OAI21_X1 g3347 (
	   .ZN (n5169),
	   .B2 (new_n7279_),
	   .B1 (new_n10076_),
	   .A (new_n10075_) );
   INV_X1 g3346 (
	   .ZN (new_n10076_),
	   .A (_net_7435) );
   NAND2_X1 g3345 (
	   .ZN (new_n10075_),
	   .A2 (new_n9722_),
	   .A1 (new_n7272_) );
   MUX2_X1 g3344 (
	   .Z (n5164),
	   .S (new_n7538_),
	   .B (_net_271),
	   .A (_net_7797) );
   CLKBUF_X1 g3343 (
	   .Z (n5159),
	   .A (_net_7793) );
   CLKBUF_X1 g3342 (
	   .Z (n5156),
	   .A (net_6428) );
   CLKBUF_X1 g3341 (
	   .Z (n5151),
	   .A (_net_7821) );
   CLKBUF_X1 g3340 (
	   .Z (n5148),
	   .A (net_6572) );
   AOI21_X1 g3339 (
	   .ZN (n5143),
	   .B2 (new_n7326_1_),
	   .B1 (new_n10068_),
	   .A (new_n10067_) );
   INV_X1 g3338 (
	   .ZN (new_n10068_),
	   .A (_net_7272) );
   NOR2_X1 g3337 (
	   .ZN (new_n10067_),
	   .A2 (n2913),
	   .A1 (new_n7325_) );
   CLKBUF_X1 g3336 (
	   .Z (n5139),
	   .A (net_6985) );
   NAND2_X1 g3335 (
	   .ZN (n5134),
	   .A2 (new_n10064_),
	   .A1 (new_n10063_) );
   AOI22_X1 g3334 (
	   .ZN (new_n10064_),
	   .B2 (net_7522),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7490) );
   AOI22_X1 g3333 (
	   .ZN (new_n10063_),
	   .B2 (_net_7426),
	   .B1 (new_n7298_),
	   .A2 (net_7458),
	   .A1 (new_n7296_) );
   AOI211_X1 g3332 (
	   .ZN (n5130),
	   .C2 (new_n7424_),
	   .C1 (new_n7182_1_),
	   .B (new_n7177_1_),
	   .A (x149) );
   CLKBUF_X1 g3331 (
	   .Z (n5126),
	   .A (net_6589) );
   CLKBUF_X1 g3330 (
	   .Z (n5121),
	   .A (net_6391) );
   NOR2_X1 g3329 (
	   .ZN (n5117),
	   .A2 (new_n7936_),
	   .A1 (new_n10058_) );
   INV_X1 g3328 (
	   .ZN (new_n10058_),
	   .A (n4304) );
   NOR3_X1 g3327 (
	   .ZN (n5112),
	   .A3 (new_n10056_1_),
	   .A2 (new_n10055_),
	   .A1 (new_n10054_) );
   INV_X1 g3326 (
	   .ZN (new_n10056_1_),
	   .A (net_6417) );
   AOI21_X1 g3325 (
	   .ZN (new_n10055_),
	   .B2 (new_n10053_),
	   .B1 (new_n7447_),
	   .A (_net_6415) );
   AND3_X1 g3324 (
	   .ZN (new_n10054_),
	   .A3 (new_n10053_),
	   .A2 (_net_6415),
	   .A1 (new_n7447_) );
   NOR2_X1 g3323 (
	   .ZN (new_n10053_),
	   .A2 (new_n10052_1_),
	   .A1 (new_n10051_) );
   INV_X1 g3322 (
	   .ZN (new_n10052_1_),
	   .A (_net_6414) );
   NAND2_X1 g3321 (
	   .ZN (new_n10051_),
	   .A2 (_net_6413),
	   .A1 (net_6412) );
   OAI221_X1 g3320 (
	   .ZN (n5107),
	   .C2 (new_n7303_),
	   .C1 (new_n9794_),
	   .B2 (new_n7306_),
	   .B1 (new_n7756_1_),
	   .A (new_n10049_) );
   AOI22_X1 g3319 (
	   .ZN (new_n10049_),
	   .B2 (_net_7416),
	   .B1 (new_n9203_),
	   .A2 (_net_7448),
	   .A1 (new_n8694_1_) );
   NAND4_X1 g3318 (
	   .ZN (n5103),
	   .A4 (new_n10047_1_),
	   .A3 (new_n10046_),
	   .A2 (new_n10045_),
	   .A1 (new_n10044_) );
   NAND4_X1 g3317 (
	   .ZN (new_n10047_1_),
	   .A4 (net_7710),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   OR2_X1 g3316 (
	   .ZN (new_n10046_),
	   .A2 (new_n7201_),
	   .A1 (new_n7365_) );
   OR2_X1 g3315 (
	   .ZN (new_n10045_),
	   .A2 (new_n7215_),
	   .A1 (new_n7362_) );
   NOR2_X1 g3314 (
	   .ZN (new_n10044_),
	   .A2 (new_n10043_),
	   .A1 (new_n10042_1_) );
   AND2_X1 g3313 (
	   .ZN (new_n10043_),
	   .A2 (net_7739),
	   .A1 (new_n7934_) );
   NAND4_X1 g3312 (
	   .ZN (new_n10042_1_),
	   .A4 (new_n10041_),
	   .A3 (new_n10040_),
	   .A2 (new_n10039_),
	   .A1 (new_n10038_) );
   NAND4_X1 g3311 (
	   .ZN (new_n10041_),
	   .A4 (_net_175),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g3310 (
	   .ZN (new_n10040_),
	   .A3 (_net_212),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g3309 (
	   .ZN (new_n10039_),
	   .A3 (net_249),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   NAND4_X1 g3308 (
	   .ZN (new_n10038_),
	   .A4 (new_n7354_1_),
	   .A3 (net_149),
	   .A2 (x1261),
	   .A1 (new_n7370_) );
   CLKBUF_X1 g3307 (
	   .Z (n5098),
	   .A (net_6399) );
   OAI21_X1 g3306 (
	   .ZN (n5094),
	   .B2 (new_n7279_),
	   .B1 (new_n10035_),
	   .A (new_n10034_) );
   INV_X1 g3305 (
	   .ZN (new_n10035_),
	   .A (_net_7433) );
   NAND2_X1 g3304 (
	   .ZN (new_n10034_),
	   .A2 (new_n7874_),
	   .A1 (new_n7272_) );
   CLKBUF_X1 g3303 (
	   .Z (n5090),
	   .A (net_7011) );
   AOI21_X1 g3302 (
	   .ZN (n5085),
	   .B2 (net_305),
	   .B1 (_net_6029),
	   .A (new_n10031_) );
   NAND3_X1 g3301 (
	   .ZN (new_n10031_),
	   .A3 (_net_6028),
	   .A2 (new_n10030_),
	   .A1 (new_n7655_) );
   INV_X1 g3300 (
	   .ZN (new_n10030_),
	   .A (net_7758) );
   OAI21_X1 g3299 (
	   .ZN (n5080),
	   .B2 (new_n7736_),
	   .B1 (new_n10028_1_),
	   .A (new_n10027_) );
   INV_X1 g3298 (
	   .ZN (new_n10028_1_),
	   .A (_net_7514) );
   NAND2_X1 g3297 (
	   .ZN (new_n10027_),
	   .A2 (new_n9502_1_),
	   .A1 (new_n7733_) );
   OAI21_X1 g3296 (
	   .ZN (n5075),
	   .B2 (new_n7736_),
	   .B1 (new_n7526_),
	   .A (new_n10025_) );
   NAND2_X1 g3295 (
	   .ZN (new_n10025_),
	   .A2 (new_n7649_1_),
	   .A1 (new_n7733_) );
   CLKBUF_X1 g3294 (
	   .Z (n5070),
	   .A (_net_7801) );
   CLKBUF_X1 g3293 (
	   .Z (n5066),
	   .A (_net_6115) );
   OAI21_X1 g3292 (
	   .ZN (n5061),
	   .B2 (new_n7736_),
	   .B1 (new_n7931_),
	   .A (new_n10021_) );
   NAND2_X1 g3291 (
	   .ZN (new_n10021_),
	   .A2 (new_n9804_),
	   .A1 (new_n7733_) );
   NOR2_X1 g3290 (
	   .ZN (n5056),
	   .A2 (new_n7334_),
	   .A1 (new_n8675_) );
   CLKBUF_X1 g3289 (
	   .Z (n5053),
	   .A (net_6970) );
   NOR2_X1 g3288 (
	   .ZN (n5048),
	   .A2 (new_n8000_),
	   .A1 (new_n7020_) );
   CLKBUF_X1 g3287 (
	   .Z (n5045),
	   .A (net_7399) );
   MUX2_X1 g3286 (
	   .Z (n5040),
	   .S (new_n6823_),
	   .B (_net_6034),
	   .A (net_7799) );
   CLKBUF_X1 g3285 (
	   .Z (n5035),
	   .A (_net_7817) );
   CLKBUF_X1 g3284 (
	   .Z (n5031),
	   .A (_net_7819) );
   NOR2_X1 g3283 (
	   .ZN (n5027),
	   .A2 (new_n6934_1_),
	   .A1 (new_n7035_) );
   CLKBUF_X1 g3282 (
	   .Z (n5023),
	   .A (net_7539) );
   AOI21_X1 g3281 (
	   .ZN (n5018),
	   .B2 (new_n10009_),
	   .B1 (_net_6693),
	   .A (new_n10010_1_) );
   OAI21_X1 g3280 (
	   .ZN (new_n10010_1_),
	   .B2 (_net_6693),
	   .B1 (new_n10009_),
	   .A (_net_5995) );
   NOR3_X1 g3279 (
	   .ZN (new_n10009_),
	   .A3 (new_n10008_),
	   .A2 (new_n7148_),
	   .A1 (new_n7228_) );
   INV_X1 g3278 (
	   .ZN (new_n10008_),
	   .A (_net_6692) );
   AOI21_X1 g3277 (
	   .ZN (n5013),
	   .B2 (new_n10006_1_),
	   .B1 (new_n10005_),
	   .A (new_n7428_) );
   INV_X1 g3276 (
	   .ZN (new_n10006_1_),
	   .A (_net_6005) );
   INV_X1 g3275 (
	   .ZN (new_n10005_),
	   .A (_net_7727) );
   CLKBUF_X1 g3274 (
	   .Z (n5008),
	   .A (net_6386) );
   CLKBUF_X1 g3273 (
	   .Z (n5005),
	   .A (net_6854) );
   CLKBUF_X1 g3272 (
	   .Z (n5001),
	   .A (net_6617) );
   CLKBUF_X1 g3271 (
	   .Z (n4996),
	   .A (_net_6065) );
   NAND3_X1 g3270 (
	   .ZN (n4992),
	   .A3 (new_n9999_),
	   .A2 (new_n9994_),
	   .A1 (new_n9985_1_) );
   AND3_X1 g3269 (
	   .ZN (new_n9999_),
	   .A3 (new_n9998_),
	   .A2 (new_n9997_1_),
	   .A1 (new_n9996_) );
   NAND2_X1 g3268 (
	   .ZN (new_n9998_),
	   .A2 (_net_7721),
	   .A1 (new_n7934_) );
   NAND4_X1 g3267 (
	   .ZN (new_n9997_1_),
	   .A4 (new_n7371_),
	   .A3 (new_n7370_),
	   .A2 (_net_6029),
	   .A1 (new_n7369_) );
   NAND2_X1 g3266 (
	   .ZN (new_n9996_),
	   .A2 (_net_115),
	   .A1 (new_n9995_) );
   INV_X1 g3265 (
	   .ZN (new_n9995_),
	   .A (new_n7374_) );
   NOR2_X1 g3264 (
	   .ZN (new_n9994_),
	   .A2 (new_n9993_),
	   .A1 (new_n9987_) );
   NAND4_X1 g3263 (
	   .ZN (new_n9993_),
	   .A4 (new_n9992_1_),
	   .A3 (new_n9991_),
	   .A2 (new_n9990_),
	   .A1 (new_n9989_) );
   NAND3_X1 g3262 (
	   .ZN (new_n9992_1_),
	   .A3 (net_194),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND4_X1 g3261 (
	   .ZN (new_n9991_),
	   .A4 (net_157),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g3260 (
	   .ZN (new_n9990_),
	   .A3 (net_231),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   NAND4_X1 g3259 (
	   .ZN (new_n9989_),
	   .A4 (new_n9988_1_),
	   .A3 (x38),
	   .A2 (new_n7381_1_),
	   .A1 (new_n7370_) );
   NAND2_X1 g3258 (
	   .ZN (new_n9988_1_),
	   .A2 (x1215),
	   .A1 (new_n7356_) );
   NOR2_X1 g3257 (
	   .ZN (new_n9987_),
	   .A2 (new_n9986_),
	   .A1 (new_n7362_) );
   INV_X1 g3256 (
	   .ZN (new_n9986_),
	   .A (_net_268) );
   NOR2_X1 g3255 (
	   .ZN (new_n9985_1_),
	   .A2 (new_n9984_),
	   .A1 (new_n9982_) );
   NOR2_X1 g3254 (
	   .ZN (new_n9984_),
	   .A2 (new_n9983_),
	   .A1 (new_n7366_) );
   INV_X1 g3253 (
	   .ZN (new_n9983_),
	   .A (_net_5985) );
   NOR2_X1 g3252 (
	   .ZN (new_n9982_),
	   .A2 (new_n9981_1_),
	   .A1 (new_n9215_1_) );
   INV_X1 g3251 (
	   .ZN (new_n9981_1_),
	   .A (_net_7692) );
   MUX2_X1 g3250 (
	   .Z (n4987),
	   .S (new_n7609_),
	   .B (_net_7571),
	   .A (new_n7216_1_) );
   CLKBUF_X1 g3249 (
	   .Z (n4983),
	   .A (net_6858) );
   CLKBUF_X1 g3248 (
	   .Z (n4979),
	   .A (net_6484) );
   NAND3_X1 g3247 (
	   .ZN (n4974),
	   .A3 (new_n9976_1_),
	   .A2 (new_n9975_),
	   .A1 (new_n9966_1_) );
   AOI22_X1 g3246 (
	   .ZN (new_n9976_1_),
	   .B2 (new_n8180_),
	   .B1 (net_7085),
	   .A2 (new_n8171_),
	   .A1 (new_n7060_) );
   AND3_X1 g3245 (
	   .ZN (new_n9975_),
	   .A3 (new_n9974_),
	   .A2 (new_n9973_),
	   .A1 (new_n9967_) );
   NAND2_X1 g3244 (
	   .ZN (new_n9974_),
	   .A2 (_net_6157),
	   .A1 (new_n7092_) );
   NAND2_X1 g3243 (
	   .ZN (new_n9973_),
	   .A2 (new_n7088_),
	   .A1 (new_n9972_) );
   NAND4_X1 g3242 (
	   .ZN (new_n9972_),
	   .A4 (new_n9971_1_),
	   .A3 (new_n9970_),
	   .A2 (new_n9969_),
	   .A1 (new_n9968_) );
   NAND3_X1 g3241 (
	   .ZN (new_n9971_1_),
	   .A3 (_net_7093),
	   .A2 (net_7073),
	   .A1 (_net_7094) );
   NAND3_X1 g3240 (
	   .ZN (new_n9970_),
	   .A3 (net_7041),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g3239 (
	   .ZN (new_n9969_),
	   .A3 (net_7009),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   NAND2_X1 g3238 (
	   .ZN (new_n9968_),
	   .A2 (net_6977),
	   .A1 (new_n7063_) );
   NAND2_X1 g3237 (
	   .ZN (new_n9967_),
	   .A2 (new_n7070_),
	   .A1 (new_n8165_) );
   AND3_X1 g3236 (
	   .ZN (new_n9966_1_),
	   .A3 (new_n9965_),
	   .A2 (new_n9964_),
	   .A1 (new_n9963_) );
   NAND4_X1 g3235 (
	   .ZN (new_n9965_),
	   .A4 (new_n7044_),
	   .A3 (net_7053),
	   .A2 (_net_7092),
	   .A1 (new_n8158_) );
   NAND4_X1 g3234 (
	   .ZN (new_n9964_),
	   .A4 (new_n7052_),
	   .A3 (_net_7092),
	   .A2 (net_6989),
	   .A1 (new_n8158_) );
   NAND4_X1 g3233 (
	   .ZN (new_n9963_),
	   .A4 (new_n7050_),
	   .A3 (net_7021),
	   .A2 (_net_7092),
	   .A1 (new_n8155_) );
   CLKBUF_X1 g3232 (
	   .Z (n4969),
	   .A (_net_7811) );
   CLKBUF_X1 g3231 (
	   .Z (n4965),
	   .A (_net_7823) );
   MUX2_X1 g3230 (
	   .Z (n4961),
	   .S (new_n7545_),
	   .B (_net_7651),
	   .A (new_n9197_) );
   CLKBUF_X1 g3229 (
	   .Z (n4957),
	   .A (net_6718) );
   MUX2_X1 g3228 (
	   .Z (n4952),
	   .S (new_n7538_),
	   .B (_net_295),
	   .A (_net_7815) );
   CLKBUF_X1 g3227 (
	   .Z (n4947),
	   .A (_net_7818) );
   CLKBUF_X1 g3226 (
	   .Z (n4944),
	   .A (net_7807) );
   CLKBUF_X1 g3225 (
	   .Z (n4940),
	   .A (_net_7812) );
   MUX2_X1 g3224 (
	   .Z (n4936),
	   .S (new_n7545_),
	   .B (_net_7659),
	   .A (new_n7022_) );
   CLKBUF_X1 g3223 (
	   .Z (n4931),
	   .A (_net_7823) );
   OAI21_X1 g3222 (
	   .ZN (n4927),
	   .B2 (new_n9338_),
	   .B1 (new_n9951_),
	   .A (new_n9949_1_) );
   NAND3_X1 g3221 (
	   .ZN (new_n9951_),
	   .A3 (new_n9950_),
	   .A2 (new_n9342_),
	   .A1 (new_n9344_) );
   NAND2_X1 g3220 (
	   .ZN (new_n9950_),
	   .A2 (_net_7782),
	   .A1 (_net_7781) );
   OAI211_X1 g3219 (
	   .ZN (new_n9949_1_),
	   .C2 (new_n9338_),
	   .C1 (new_n9341_),
	   .B (_net_7782),
	   .A (new_n9342_) );
   XNOR2_X1 g3218 (
	   .ZN (n4922),
	   .B (new_n8395_),
	   .A (new_n8393_) );
   MUX2_X1 g3217 (
	   .Z (n4917),
	   .S (new_n7437_1_),
	   .B (_net_6011),
	   .A (_net_7814) );
   CLKBUF_X1 g3216 (
	   .Z (n4913),
	   .A (net_6573) );
   NOR2_X1 g3215 (
	   .ZN (n4908),
	   .A2 (new_n8387_1_),
	   .A1 (new_n9927_) );
   CLKBUF_X1 g3214 (
	   .Z (n4904),
	   .A (net_7001) );
   CLKBUF_X1 g3213 (
	   .Z (n4899),
	   .A (_net_6143) );
   CLKBUF_X1 g3212 (
	   .Z (n4895),
	   .A (net_7154) );
   CLKBUF_X1 g3211 (
	   .Z (n4890),
	   .A (_net_7801) );
   OAI221_X1 g3210 (
	   .ZN (n4886),
	   .C2 (new_n7306_),
	   .C1 (new_n9939_1_),
	   .B2 (new_n7303_),
	   .B1 (new_n6937_),
	   .A (new_n9938_) );
   INV_X1 g3209 (
	   .ZN (new_n9939_1_),
	   .A (_net_7506) );
   AOI22_X1 g3208 (
	   .ZN (new_n9938_),
	   .B2 (_net_7410),
	   .B1 (new_n9203_),
	   .A2 (_net_7442),
	   .A1 (new_n8694_1_) );
   CLKBUF_X1 g3207 (
	   .Z (n4881),
	   .A (net_6384) );
   OAI21_X1 g3206 (
	   .ZN (n4877),
	   .B2 (new_n9935_1_),
	   .B1 (new_n9934_),
	   .A (new_n6963_) );
   INV_X1 g3205 (
	   .ZN (new_n9935_1_),
	   .A (new_n9303_) );
   NOR2_X1 g3204 (
	   .ZN (new_n9934_),
	   .A2 (_net_6406),
	   .A1 (new_n9933_) );
   NOR2_X1 g3203 (
	   .ZN (new_n9933_),
	   .A2 (new_n9683_1_),
	   .A1 (new_n8188_1_) );
   MUX2_X1 g3202 (
	   .Z (n4872),
	   .S (new_n7538_),
	   .B (_net_284),
	   .A (net_7807) );
   CLKBUF_X1 g3201 (
	   .Z (n4867),
	   .A (_net_7819) );
   CLKBUF_X1 g3200 (
	   .Z (n4862),
	   .A (_net_6402) );
   NOR2_X1 g3199 (
	   .ZN (n4857),
	   .A2 (new_n9928_),
	   .A1 (new_n9927_) );
   INV_X1 g3198 (
	   .ZN (new_n9928_),
	   .A (new_n6820_) );
   NAND3_X1 g3197 (
	   .ZN (new_n9927_),
	   .A3 (new_n7389_),
	   .A2 (x1231),
	   .A1 (new_n7183_) );
   CLKBUF_X1 g3196 (
	   .Z (n4853),
	   .A (net_6875) );
   CLKBUF_X1 g3195 (
	   .Z (n4848),
	   .A (_net_6074) );
   MUX2_X1 g3194 (
	   .Z (n4843),
	   .S (new_n7437_1_),
	   .B (_net_6019),
	   .A (_net_7819) );
   CLKBUF_X1 g3193 (
	   .Z (n4838),
	   .A (_net_7814) );
   CLKBUF_X1 g3192 (
	   .Z (n4834),
	   .A (_net_7820) );
   OAI211_X1 g3191 (
	   .ZN (n4831),
	   .C2 (new_n7366_),
	   .C1 (new_n6861_),
	   .B (new_n9920_),
	   .A (new_n9919_) );
   NAND4_X1 g3190 (
	   .ZN (new_n9920_),
	   .A4 (_net_7717),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   NOR3_X1 g3189 (
	   .ZN (new_n9919_),
	   .A3 (new_n9918_1_),
	   .A2 (new_n9917_),
	   .A1 (new_n9916_) );
   AND3_X1 g3188 (
	   .ZN (new_n9918_1_),
	   .A3 (new_n7382_),
	   .A2 (net_256),
	   .A1 (new_n7380_) );
   NOR2_X1 g3187 (
	   .ZN (new_n9917_),
	   .A2 (new_n7891_),
	   .A1 (new_n7378_) );
   OAI22_X1 g3186 (
	   .ZN (new_n9916_),
	   .B2 (new_n9915_),
	   .B1 (new_n7938_),
	   .A2 (new_n9914_1_),
	   .A1 (new_n7936_) );
   INV_X1 g3185 (
	   .ZN (new_n9915_),
	   .A (net_182) );
   INV_X1 g3184 (
	   .ZN (new_n9914_1_),
	   .A (net_219) );
   CLKBUF_X1 g3183 (
	   .Z (n4827),
	   .A (net_6567) );
   NOR2_X1 g3182 (
	   .ZN (n4822),
	   .A2 (new_n7494_),
	   .A1 (new_n8675_) );
   MUX2_X1 g3181 (
	   .Z (n4818),
	   .S (new_n7504_),
	   .B (_net_7624),
	   .A (new_n9910_) );
   OAI21_X1 g3180 (
	   .ZN (new_n9910_),
	   .B2 (new_n9909_),
	   .B1 (new_n7019_),
	   .A (new_n9908_) );
   INV_X1 g3179 (
	   .ZN (new_n9909_),
	   .A (net_7544) );
   AOI22_X1 g3178 (
	   .ZN (new_n9908_),
	   .B2 (net_374),
	   .B1 (_net_292),
	   .A2 (_net_291),
	   .A1 (net_376) );
   CLKBUF_X1 g3177 (
	   .Z (n4814),
	   .A (net_7128) );
   MUX2_X1 g3176 (
	   .Z (n4809),
	   .S (new_n7545_),
	   .B (_net_7655),
	   .A (new_n9509_) );
   CLKBUF_X1 g3175 (
	   .Z (n4805),
	   .A (net_7014) );
   OAI21_X1 g3174 (
	   .ZN (n4800),
	   .B2 (new_n7279_),
	   .B1 (new_n9903_),
	   .A (new_n9902_1_) );
   INV_X1 g3173 (
	   .ZN (new_n9903_),
	   .A (_net_7452) );
   NAND2_X1 g3172 (
	   .ZN (new_n9902_1_),
	   .A2 (new_n9901_),
	   .A1 (new_n7272_) );
   OAI22_X1 g3171 (
	   .ZN (new_n9901_),
	   .B2 (new_n6901_),
	   .B1 (new_n9900_),
	   .A2 (new_n7962_1_),
	   .A1 (new_n7034_) );
   INV_X1 g3170 (
	   .ZN (new_n9900_),
	   .A (net_365) );
   CLKBUF_X1 g3169 (
	   .Z (n4795),
	   .A (_net_7803) );
   CLKBUF_X1 g3168 (
	   .Z (n4791),
	   .A (net_7799) );
   MUX2_X1 g3167 (
	   .Z (n4787),
	   .S (new_n7609_),
	   .B (_net_7559),
	   .A (new_n9509_) );
   CLKBUF_X1 g3166 (
	   .Z (n4782),
	   .A (_net_6156) );
   CLKBUF_X1 g3165 (
	   .Z (n4778),
	   .A (net_6449) );
   CLKBUF_X1 g3164 (
	   .Z (n4774),
	   .A (net_7545) );
   NOR2_X1 g3163 (
	   .ZN (n4769),
	   .A2 (new_n7274_),
	   .A1 (new_n8543_) );
   CLKBUF_X1 g3162 (
	   .Z (n4765),
	   .A (net_137) );
   MUX2_X1 g3161 (
	   .Z (n4760),
	   .S (new_n7285_),
	   .B (_net_7706),
	   .A (_net_7808) );
   CLKBUF_X1 g3160 (
	   .Z (n4755),
	   .A (_net_6153) );
   CLKBUF_X1 g3159 (
	   .Z (n4750),
	   .A (_net_6138) );
   CLKBUF_X1 g3158 (
	   .Z (n4745),
	   .A (net_7807) );
   CLKBUF_X1 g3157 (
	   .Z (n4742),
	   .A (net_6735) );
   AOI21_X1 g3156 (
	   .ZN (n4737),
	   .B2 (new_n6945_),
	   .B1 (_net_7382),
	   .A (new_n9885_1_) );
   OAI21_X1 g3155 (
	   .ZN (new_n9885_1_),
	   .B2 (_net_7382),
	   .B1 (new_n6945_),
	   .A (_net_267) );
   OAI21_X1 g3154 (
	   .ZN (n4732),
	   .B2 (new_n7258_),
	   .B1 (new_n7311_),
	   .A (new_n9883_) );
   NAND2_X1 g3153 (
	   .ZN (new_n9883_),
	   .A2 (new_n9002_),
	   .A1 (new_n7252_1_) );
   OAI21_X1 g3152 (
	   .ZN (n4727),
	   .B2 (new_n7285_),
	   .B1 (new_n8091_),
	   .A (new_n9881_) );
   NAND2_X1 g3151 (
	   .ZN (new_n9881_),
	   .A2 (_net_7692),
	   .A1 (new_n7285_) );
   CLKBUF_X1 g3150 (
	   .Z (n4722),
	   .A (_net_6095) );
   CLKBUF_X1 g3149 (
	   .Z (n4717),
	   .A (_net_7817) );
   CLKBUF_X1 g3148 (
	   .Z (n4713),
	   .A (net_7142) );
   NAND3_X1 g3147 (
	   .ZN (n4708),
	   .A3 (new_n9876_),
	   .A2 (new_n9872_),
	   .A1 (new_n9868_) );
   AND3_X1 g3146 (
	   .ZN (new_n9876_),
	   .A3 (new_n9875_1_),
	   .A2 (new_n9874_),
	   .A1 (new_n9873_) );
   NAND2_X1 g3145 (
	   .ZN (new_n9875_1_),
	   .A2 (_net_6073),
	   .A1 (new_n6813_1_) );
   NAND2_X1 g3144 (
	   .ZN (new_n9874_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n9238_1_) );
   NAND2_X1 g3143 (
	   .ZN (new_n9873_),
	   .A2 (new_n7166_),
	   .A1 (new_n8079_) );
   AOI22_X1 g3142 (
	   .ZN (new_n9872_),
	   .B2 (net_6541),
	   .B1 (new_n6779_1_),
	   .A2 (new_n6784_),
	   .A1 (new_n9871_1_) );
   NAND2_X1 g3141 (
	   .ZN (new_n9871_1_),
	   .A2 (new_n9870_),
	   .A1 (new_n9869_) );
   AOI22_X1 g3140 (
	   .ZN (new_n9870_),
	   .B2 (net_6429),
	   .B1 (new_n6785_),
	   .A2 (net_6461),
	   .A1 (new_n6766_) );
   AOI22_X1 g3139 (
	   .ZN (new_n9869_),
	   .B2 (net_6525),
	   .B1 (new_n8139_),
	   .A2 (new_n6774_1_),
	   .A1 (net_6493) );
   AND3_X1 g3138 (
	   .ZN (new_n9868_),
	   .A3 (new_n9867_1_),
	   .A2 (new_n9866_),
	   .A1 (new_n9865_) );
   NAND4_X1 g3137 (
	   .ZN (new_n9867_1_),
	   .A4 (new_n6775_),
	   .A3 (_net_6552),
	   .A2 (net_6509),
	   .A1 (new_n6772_) );
   NAND4_X1 g3136 (
	   .ZN (new_n9866_),
	   .A4 (new_n6770_1_),
	   .A3 (net_6445),
	   .A2 (_net_6552),
	   .A1 (new_n6772_) );
   NAND4_X1 g3135 (
	   .ZN (new_n9865_),
	   .A4 (new_n6767_),
	   .A3 (_net_6552),
	   .A2 (net_6477),
	   .A1 (new_n6764_) );
   INV_X1 g3134 (
	   .ZN (n4703),
	   .A (new_n6780_) );
   CLKBUF_X1 g3133 (
	   .Z (n4699),
	   .A (net_6993) );
   NOR2_X1 g3132 (
	   .ZN (n4694),
	   .A2 (new_n6900_),
	   .A1 (new_n8543_) );
   AND2_X1 g3131 (
	   .ZN (n4690),
	   .A2 (net_338),
	   .A1 (new_n7102_1_) );
   CLKBUF_X1 g3130 (
	   .Z (n4686),
	   .A (net_6393) );
   CLKBUF_X1 g3129 (
	   .Z (n4681),
	   .A (x1564) );
   NAND3_X1 g3128 (
	   .ZN (n4678),
	   .A3 (new_n9857_),
	   .A2 (new_n9856_),
	   .A1 (new_n9848_) );
   NAND4_X1 g3127 (
	   .ZN (new_n9857_),
	   .A4 (_net_7693),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR3_X1 g3126 (
	   .ZN (new_n9856_),
	   .A3 (new_n9855_),
	   .A2 (new_n9851_),
	   .A1 (new_n9849_1_) );
   NAND3_X1 g3125 (
	   .ZN (new_n9855_),
	   .A3 (new_n9854_),
	   .A2 (new_n9853_1_),
	   .A1 (new_n9852_) );
   NAND4_X1 g3124 (
	   .ZN (new_n9854_),
	   .A4 (net_158),
	   .A3 (x1231),
	   .A2 (new_n7394_),
	   .A1 (new_n7392_) );
   NAND3_X1 g3123 (
	   .ZN (new_n9853_1_),
	   .A3 (net_195),
	   .A2 (new_n7388_),
	   .A1 (new_n7386_1_) );
   NAND3_X1 g3122 (
	   .ZN (new_n9852_),
	   .A3 (net_232),
	   .A2 (new_n7382_),
	   .A1 (new_n7380_) );
   OAI22_X1 g3121 (
	   .ZN (new_n9851_),
	   .B2 (new_n7378_),
	   .B1 (new_n8873_1_),
	   .A2 (new_n9850_),
	   .A1 (new_n7374_) );
   INV_X1 g3120 (
	   .ZN (new_n9850_),
	   .A (_net_116) );
   AND4_X1 g3119 (
	   .ZN (new_n9849_1_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7369_),
	   .A1 (_net_6030) );
   NOR2_X1 g3118 (
	   .ZN (new_n9848_),
	   .A2 (new_n9847_),
	   .A1 (new_n9846_) );
   NOR2_X1 g3117 (
	   .ZN (new_n9847_),
	   .A2 (new_n6799_),
	   .A1 (new_n7366_) );
   NOR2_X1 g3116 (
	   .ZN (new_n9846_),
	   .A2 (new_n7105_),
	   .A1 (new_n7362_) );
   NOR4_X1 g3115 (
	   .ZN (n4673),
	   .A4 (_net_6410),
	   .A3 (new_n8183_1_),
	   .A2 (new_n8187_),
	   .A1 (new_n9844_1_) );
   NAND4_X1 g3114 (
	   .ZN (new_n9844_1_),
	   .A4 (_net_6407),
	   .A3 (_net_6404),
	   .A2 (new_n9683_1_),
	   .A1 (new_n9682_) );
   CLKBUF_X1 g3113 (
	   .Z (n4669),
	   .A (net_6581) );
   CLKBUF_X1 g3112 (
	   .Z (n4665),
	   .A (net_6736) );
   CLKBUF_X1 g3111 (
	   .Z (n4660),
	   .A (_net_7795) );
   OAI21_X1 g3110 (
	   .ZN (n4656),
	   .B2 (new_n7258_),
	   .B1 (new_n9839_),
	   .A (new_n9838_) );
   INV_X1 g3109 (
	   .ZN (new_n9839_),
	   .A (_net_7288) );
   NAND2_X1 g3108 (
	   .ZN (new_n9838_),
	   .A2 (new_n8292_),
	   .A1 (new_n7252_1_) );
   CLKBUF_X1 g3107 (
	   .Z (n4651),
	   .A (_net_6171) );
   OAI21_X1 g3106 (
	   .ZN (n4646),
	   .B2 (new_n6957_1_),
	   .B1 (new_n9835_),
	   .A (new_n9834_) );
   INV_X1 g3105 (
	   .ZN (new_n9835_),
	   .A (_net_7269) );
   NAND2_X1 g3104 (
	   .ZN (new_n9834_),
	   .A2 (new_n9707_),
	   .A1 (new_n6949_) );
   OAI21_X1 g3103 (
	   .ZN (n4641),
	   .B2 (new_n9469_),
	   .B1 (new_n9832_),
	   .A (new_n9831_) );
   INV_X1 g3102 (
	   .ZN (new_n9832_),
	   .A (_net_6064) );
   NAND2_X1 g3101 (
	   .ZN (new_n9831_),
	   .A2 (new_n7166_),
	   .A1 (new_n9830_) );
   NAND2_X1 g3100 (
	   .ZN (new_n9830_),
	   .A2 (new_n9829_),
	   .A1 (new_n9828_1_) );
   AOI22_X1 g3099 (
	   .ZN (new_n9829_),
	   .B2 (net_6424),
	   .B1 (new_n6770_1_),
	   .A2 (net_6456),
	   .A1 (new_n6766_) );
   AOI22_X1 g3098 (
	   .ZN (new_n9828_1_),
	   .B2 (net_6520),
	   .B1 (new_n8139_),
	   .A2 (new_n6774_1_),
	   .A1 (net_6488) );
   NAND2_X1 g3097 (
	   .ZN (n4636),
	   .A2 (new_n9826_),
	   .A1 (new_n9825_) );
   AOI22_X1 g3096 (
	   .ZN (new_n9826_),
	   .B2 (_net_7575),
	   .B1 (new_n6755_),
	   .A2 (net_7607),
	   .A1 (new_n6743_) );
   AOI22_X1 g3095 (
	   .ZN (new_n9825_),
	   .B2 (net_7639),
	   .B1 (new_n8009_),
	   .A2 (new_n7970_1_),
	   .A1 (net_7671) );
   CLKBUF_X1 g3094 (
	   .Z (n4631),
	   .A (_net_7821) );
   OAI21_X1 g3093 (
	   .ZN (n4627),
	   .B2 (new_n7111_1_),
	   .B1 (new_n9822_),
	   .A (new_n9821_) );
   INV_X1 g3092 (
	   .ZN (new_n9822_),
	   .A (_net_7346) );
   NAND2_X1 g3091 (
	   .ZN (new_n9821_),
	   .A2 (new_n8780_1_),
	   .A1 (new_n7101_) );
   CLKBUF_X1 g3090 (
	   .Z (n4622),
	   .A (_net_6097) );
   CLKBUF_X1 g3089 (
	   .Z (n4617),
	   .A (net_7807) );
   CLKBUF_X1 g3088 (
	   .Z (n4613),
	   .A (_net_7811) );
   MUX2_X1 g3087 (
	   .Z (n4609),
	   .S (new_n7029_),
	   .B (_net_7586),
	   .A (new_n8114_) );
   CLKBUF_X1 g3086 (
	   .Z (n4604),
	   .A (_net_7805) );
   CLKBUF_X1 g3085 (
	   .Z (n4600),
	   .A (_net_7801) );
   OAI21_X1 g3084 (
	   .ZN (n4596),
	   .B2 (new_n7652_),
	   .B1 (new_n9813_),
	   .A (new_n9812_) );
   INV_X1 g3083 (
	   .ZN (new_n9813_),
	   .A (_net_7413) );
   NAND2_X1 g3082 (
	   .ZN (new_n9812_),
	   .A2 (new_n8679_),
	   .A1 (new_n7646_) );
   AOI21_X1 g3081 (
	   .ZN (n4591),
	   .B2 (new_n9590_),
	   .B1 (_net_7233),
	   .A (new_n9810_) );
   OAI21_X1 g3080 (
	   .ZN (new_n9810_),
	   .B2 (_net_7233),
	   .B1 (new_n9590_),
	   .A (_net_6039) );
   AND2_X1 g3079 (
	   .ZN (n4586),
	   .A2 (_net_6296),
	   .A1 (new_n9520_1_) );
   CLKBUF_X1 g3078 (
	   .Z (n4581),
	   .A (_net_7812) );
   CLKBUF_X1 g3077 (
	   .Z (n4577),
	   .A (_net_6109) );
   OAI21_X1 g3076 (
	   .ZN (n4572),
	   .B2 (new_n6907_),
	   .B1 (new_n7930_),
	   .A (new_n9805_1_) );
   NAND2_X1 g3075 (
	   .ZN (new_n9805_1_),
	   .A2 (new_n9804_),
	   .A1 (new_n6897_) );
   OAI221_X1 g3074 (
	   .ZN (new_n9804_),
	   .C2 (new_n6901_),
	   .C1 (new_n7274_),
	   .B2 (new_n8678_),
	   .B1 (new_n6902_1_),
	   .A (new_n9803_) );
   NAND2_X1 g3073 (
	   .ZN (new_n9803_),
	   .A2 (net_7395),
	   .A1 (new_n6889_) );
   CLKBUF_X1 g3072 (
	   .Z (n4567),
	   .A (net_131) );
   CLKBUF_X1 g3071 (
	   .Z (n4562),
	   .A (_net_7796) );
   CLKBUF_X1 g3070 (
	   .Z (n4558),
	   .A (_net_7809) );
   OAI21_X1 g3069 (
	   .ZN (n4553),
	   .B2 (new_n7692_),
	   .B1 (new_n9798_),
	   .A (new_n9797_) );
   INV_X1 g3068 (
	   .ZN (new_n9798_),
	   .A (_net_6165) );
   NAND2_X1 g3067 (
	   .ZN (new_n9797_),
	   .A2 (new_n7690_),
	   .A1 (new_n7698_) );
   CLKBUF_X1 g3066 (
	   .Z (n4548),
	   .A (_net_7794) );
   OAI21_X1 g3065 (
	   .ZN (n4544),
	   .B2 (new_n6907_),
	   .B1 (new_n9794_),
	   .A (new_n9793_) );
   INV_X1 g3064 (
	   .ZN (new_n9794_),
	   .A (_net_7480) );
   NAND2_X1 g3063 (
	   .ZN (new_n9793_),
	   .A2 (new_n7754_),
	   .A1 (new_n6897_) );
   NAND3_X1 g3062 (
	   .ZN (n4539),
	   .A3 (new_n9791_),
	   .A2 (new_n9790_),
	   .A1 (new_n9776_) );
   AOI22_X1 g3061 (
	   .ZN (new_n9791_),
	   .B2 (new_n7844_),
	   .B1 (net_7215),
	   .A2 (new_n7837_),
	   .A1 (new_n8022_) );
   AND3_X1 g3060 (
	   .ZN (new_n9790_),
	   .A3 (new_n9789_),
	   .A2 (new_n9788_),
	   .A1 (new_n9782_) );
   NAND2_X1 g3059 (
	   .ZN (new_n9789_),
	   .A2 (_net_6172),
	   .A1 (new_n7694_) );
   NAND2_X1 g3058 (
	   .ZN (new_n9788_),
	   .A2 (new_n7701_),
	   .A1 (new_n9787_1_) );
   NAND4_X1 g3057 (
	   .ZN (new_n9787_1_),
	   .A4 (new_n9786_),
	   .A3 (new_n9785_),
	   .A2 (new_n9784_),
	   .A1 (new_n9783_1_) );
   NAND3_X1 g3056 (
	   .ZN (new_n9786_),
	   .A3 (_net_7228),
	   .A2 (_net_7229),
	   .A1 (net_7201) );
   NAND3_X1 g3055 (
	   .ZN (new_n9785_),
	   .A3 (net_7169),
	   .A2 (_net_7229),
	   .A1 (new_n7823_) );
   NAND3_X1 g3054 (
	   .ZN (new_n9784_),
	   .A3 (net_7137),
	   .A2 (_net_7228),
	   .A1 (new_n7821_) );
   NAND2_X1 g3053 (
	   .ZN (new_n9783_1_),
	   .A2 (net_7105),
	   .A1 (new_n7819_) );
   NAND2_X1 g3052 (
	   .ZN (new_n9782_),
	   .A2 (new_n7690_),
	   .A1 (new_n9781_) );
   NAND4_X1 g3051 (
	   .ZN (new_n9781_),
	   .A4 (new_n9780_),
	   .A3 (new_n9779_),
	   .A2 (new_n9778_1_),
	   .A1 (new_n9777_) );
   NAND3_X1 g3050 (
	   .ZN (new_n9780_),
	   .A3 (_net_7228),
	   .A2 (net_7203),
	   .A1 (_net_7229) );
   NAND3_X1 g3049 (
	   .ZN (new_n9779_),
	   .A3 (net_7171),
	   .A2 (_net_7229),
	   .A1 (new_n7823_) );
   NAND3_X1 g3048 (
	   .ZN (new_n9778_1_),
	   .A3 (_net_7228),
	   .A2 (net_7139),
	   .A1 (new_n7821_) );
   NAND2_X1 g3047 (
	   .ZN (new_n9777_),
	   .A2 (net_7107),
	   .A1 (new_n7819_) );
   AND3_X1 g3046 (
	   .ZN (new_n9776_),
	   .A3 (new_n9775_),
	   .A2 (new_n9774_),
	   .A1 (new_n9773_1_) );
   NAND4_X1 g3045 (
	   .ZN (new_n9775_),
	   .A4 (new_n7678_),
	   .A3 (net_7183),
	   .A2 (_net_7227),
	   .A1 (new_n7816_) );
   NAND4_X1 g3044 (
	   .ZN (new_n9774_),
	   .A4 (new_n7683_),
	   .A3 (_net_7227),
	   .A2 (net_7119),
	   .A1 (new_n7816_) );
   NAND4_X1 g3043 (
	   .ZN (new_n9773_1_),
	   .A4 (new_n7681_1_),
	   .A3 (net_7151),
	   .A2 (_net_7227),
	   .A1 (new_n7813_) );
   AND2_X1 g3042 (
	   .ZN (n4534),
	   .A2 (_net_6194),
	   .A1 (new_n9520_1_) );
   AND2_X1 g3041 (
	   .ZN (n4529),
	   .A2 (_net_6188),
	   .A1 (new_n9520_1_) );
   CLKBUF_X1 g3040 (
	   .Z (n4524),
	   .A (_net_7801) );
   NAND2_X1 g3039 (
	   .ZN (n4520),
	   .A2 (new_n9768_1_),
	   .A1 (new_n9767_) );
   AOI22_X1 g3038 (
	   .ZN (new_n9768_1_),
	   .B2 (new_n6751_),
	   .B1 (_net_7568),
	   .A2 (_net_7664),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g3037 (
	   .ZN (new_n9767_),
	   .B2 (_net_7600),
	   .B1 (new_n7350_),
	   .A2 (new_n6746_1_),
	   .A1 (_net_7632) );
   NAND3_X1 g3036 (
	   .ZN (n4515),
	   .A3 (new_n9765_),
	   .A2 (new_n9764_),
	   .A1 (new_n9760_) );
   AOI22_X1 g3035 (
	   .ZN (new_n9765_),
	   .B2 (new_n7844_),
	   .B1 (net_7216),
	   .A2 (new_n7837_),
	   .A1 (new_n8547_) );
   AND3_X1 g3034 (
	   .ZN (new_n9764_),
	   .A3 (new_n9763_1_),
	   .A2 (new_n9762_),
	   .A1 (new_n9761_) );
   NAND2_X1 g3033 (
	   .ZN (new_n9763_1_),
	   .A2 (_net_6173),
	   .A1 (new_n7694_) );
   NAND2_X1 g3032 (
	   .ZN (new_n9762_),
	   .A2 (new_n7701_),
	   .A1 (new_n9057_1_) );
   NAND2_X1 g3031 (
	   .ZN (new_n9761_),
	   .A2 (new_n7690_),
	   .A1 (new_n8376_) );
   AND3_X1 g3030 (
	   .ZN (new_n9760_),
	   .A3 (new_n9759_),
	   .A2 (new_n9758_1_),
	   .A1 (new_n9757_) );
   NAND4_X1 g3029 (
	   .ZN (new_n9759_),
	   .A4 (new_n7678_),
	   .A3 (_net_7227),
	   .A2 (net_7184),
	   .A1 (new_n7816_) );
   NAND4_X1 g3028 (
	   .ZN (new_n9758_1_),
	   .A4 (new_n7683_),
	   .A3 (_net_7227),
	   .A2 (net_7120),
	   .A1 (new_n7816_) );
   NAND4_X1 g3027 (
	   .ZN (new_n9757_),
	   .A4 (new_n7681_1_),
	   .A3 (net_7152),
	   .A2 (_net_7227),
	   .A1 (new_n7813_) );
   OAI21_X1 g3026 (
	   .ZN (n4510),
	   .B2 (new_n6907_),
	   .B1 (new_n9205_),
	   .A (new_n9755_) );
   NAND2_X1 g3025 (
	   .ZN (new_n9755_),
	   .A2 (new_n8859_),
	   .A1 (new_n6897_) );
   CLKBUF_X1 g3024 (
	   .Z (n4505),
	   .A (_net_7808) );
   NOR2_X1 g3023 (
	   .ZN (n4501),
	   .A2 (net_153),
	   .A1 (new_n9752_) );
   INV_X1 g3022 (
	   .ZN (new_n9752_),
	   .A (_net_7768) );
   CLKBUF_X1 g3021 (
	   .Z (n4496),
	   .A (net_386) );
   MUX2_X1 g3020 (
	   .Z (n4491),
	   .S (new_n7437_1_),
	   .B (_net_6018),
	   .A (_net_7818) );
   CLKBUF_X1 g3019 (
	   .Z (n4487),
	   .A (net_7129) );
   NAND4_X1 g3018 (
	   .ZN (n4482),
	   .A4 (new_n9747_),
	   .A3 (new_n9743_),
	   .A2 (new_n9742_1_),
	   .A1 (new_n9741_) );
   NAND2_X1 g3017 (
	   .ZN (new_n9747_),
	   .A2 (new_n7060_),
	   .A1 (new_n9746_1_) );
   NAND2_X1 g3016 (
	   .ZN (new_n9746_1_),
	   .A2 (new_n9745_),
	   .A1 (new_n9744_) );
   AOI22_X1 g3015 (
	   .ZN (new_n9745_),
	   .B2 (net_6964),
	   .B1 (new_n7052_),
	   .A2 (net_6996),
	   .A1 (new_n7049_1_) );
   AOI22_X1 g3014 (
	   .ZN (new_n9744_),
	   .B2 (net_7060),
	   .B1 (new_n7046_),
	   .A2 (new_n7043_),
	   .A1 (net_7028) );
   NAND2_X1 g3013 (
	   .ZN (new_n9743_),
	   .A2 (new_n8656_),
	   .A1 (new_n7073_) );
   NAND2_X1 g3012 (
	   .ZN (new_n9742_1_),
	   .A2 (new_n7070_),
	   .A1 (new_n7054_) );
   AOI22_X1 g3011 (
	   .ZN (new_n9741_),
	   .B2 (new_n7092_),
	   .B1 (_net_6148),
	   .A2 (new_n7089_1_),
	   .A1 (new_n7065_) );
   CLKBUF_X1 g3010 (
	   .Z (n4478),
	   .A (net_6448) );
   CLKBUF_X1 g3009 (
	   .Z (n4473),
	   .A (_net_7797) );
   CLKBUF_X1 g3008 (
	   .Z (n4469),
	   .A (_net_6147) );
   OAI21_X1 g3007 (
	   .ZN (n4464),
	   .B2 (new_n7225_),
	   .B1 (new_n9736_),
	   .A (new_n9735_) );
   INV_X1 g3006 (
	   .ZN (new_n9736_),
	   .A (_net_7323) );
   NAND2_X1 g3005 (
	   .ZN (new_n9735_),
	   .A2 (new_n7108_),
	   .A1 (new_n7222_) );
   NAND2_X1 g3004 (
	   .ZN (n4459),
	   .A2 (n4304),
	   .A1 (new_n7422_1_) );
   OAI221_X1 g3003 (
	   .ZN (n4456),
	   .C2 (new_n7936_),
	   .C1 (new_n9732_),
	   .B2 (new_n7366_),
	   .B1 (new_n9391_),
	   .A (new_n9731_) );
   INV_X1 g3002 (
	   .ZN (new_n9732_),
	   .A (net_223) );
   AOI22_X1 g3001 (
	   .ZN (new_n9731_),
	   .B2 (net_186),
	   .B1 (new_n9730_),
	   .A2 (new_n9729_1_),
	   .A1 (net_260) );
   INV_X1 g3000 (
	   .ZN (new_n9730_),
	   .A (new_n7938_) );
   INV_X1 g2999 (
	   .ZN (new_n9729_1_),
	   .A (new_n7369_) );
   AND2_X1 g2998 (
	   .ZN (n4451),
	   .A2 (net_342),
	   .A1 (new_n7102_1_) );
   CLKBUF_X1 g2997 (
	   .Z (n4448),
	   .A (net_6886) );
   AND2_X1 g2996 (
	   .ZN (n4443),
	   .A2 (_net_6205),
	   .A1 (new_n9520_1_) );
   OAI21_X1 g2995 (
	   .ZN (n4438),
	   .B2 (new_n7652_),
	   .B1 (new_n9724_1_),
	   .A (new_n9723_) );
   INV_X1 g2994 (
	   .ZN (new_n9724_1_),
	   .A (_net_7403) );
   NAND2_X1 g2993 (
	   .ZN (new_n9723_),
	   .A2 (new_n9722_),
	   .A1 (new_n7646_) );
   OAI21_X1 g2992 (
	   .ZN (new_n9722_),
	   .B2 (new_n9721_),
	   .B1 (new_n7034_),
	   .A (new_n9720_) );
   INV_X1 g2991 (
	   .ZN (new_n9721_),
	   .A (net_7387) );
   AOI22_X1 g2990 (
	   .ZN (new_n9720_),
	   .B2 (net_348),
	   .B1 (_net_281),
	   .A2 (net_350),
	   .A1 (_net_280) );
   OAI21_X1 g2989 (
	   .ZN (n4433),
	   .B2 (new_n7225_),
	   .B1 (new_n9718_),
	   .A (new_n9717_) );
   INV_X1 g2988 (
	   .ZN (new_n9718_),
	   .A (_net_7332) );
   NAND2_X1 g2987 (
	   .ZN (new_n9717_),
	   .A2 (new_n7335_1_),
	   .A1 (new_n7222_) );
   NOR2_X1 g2986 (
	   .ZN (n4428),
	   .A2 (new_n7493_),
	   .A1 (new_n8675_) );
   MUX2_X1 g2985 (
	   .Z (n4424),
	   .S (new_n6823_),
	   .B (_net_6045),
	   .A (net_7807) );
   CLKBUF_X1 g2984 (
	   .Z (n4419),
	   .A (_net_6151) );
   MUX2_X1 g2983 (
	   .Z (n4414),
	   .S (new_n7285_),
	   .B (_net_7718),
	   .A (_net_7820) );
   CLKBUF_X1 g2982 (
	   .Z (n4410),
	   .A (net_7111) );
   CLKBUF_X1 g2981 (
	   .Z (n4401),
	   .A (net_7162) );
   CLKBUF_X1 g2980 (
	   .Z (n4397),
	   .A (net_6564) );
   OAI21_X1 g2979 (
	   .ZN (n4392),
	   .B2 (new_n7258_),
	   .B1 (new_n6915_1_),
	   .A (new_n9708_) );
   NAND2_X1 g2978 (
	   .ZN (new_n9708_),
	   .A2 (new_n9707_),
	   .A1 (new_n7252_1_) );
   OAI22_X1 g2977 (
	   .ZN (new_n9707_),
	   .B2 (new_n7106_),
	   .B1 (new_n7602_),
	   .A2 (new_n8132_),
	   .A1 (new_n6951_) );
   CLKBUF_X1 g2976 (
	   .Z (n4388),
	   .A (net_6431) );
   CLKBUF_X1 g2975 (
	   .Z (n4384),
	   .A (net_6974) );
   AOI21_X1 g2974 (
	   .ZN (n4379),
	   .B2 (new_n7326_1_),
	   .B1 (new_n9703_),
	   .A (new_n9702_) );
   INV_X1 g2973 (
	   .ZN (new_n9703_),
	   .A (_net_7278) );
   NOR2_X1 g2972 (
	   .ZN (new_n9702_),
	   .A2 (n576),
	   .A1 (new_n7325_) );
   CLKBUF_X1 g2971 (
	   .Z (n4374),
	   .A (_net_7818) );
   CLKBUF_X1 g2970 (
	   .Z (n4370),
	   .A (_net_7811) );
   CLKBUF_X1 g2969 (
	   .Z (n4365),
	   .A (_net_7797) );
   CLKBUF_X1 g2968 (
	   .Z (n4362),
	   .A (net_6863) );
   MUX2_X1 g2967 (
	   .Z (n4357),
	   .S (new_n7437_1_),
	   .B (_net_6009),
	   .A (_net_7812) );
   NOR2_X1 g2966 (
	   .ZN (n4352),
	   .A2 (new_n8000_),
	   .A1 (new_n7020_) );
   OAI21_X1 g2965 (
	   .ZN (n4348),
	   .B2 (new_n7736_),
	   .B1 (new_n9694_),
	   .A (new_n9693_) );
   INV_X1 g2964 (
	   .ZN (new_n9694_),
	   .A (_net_7505) );
   NAND2_X1 g2963 (
	   .ZN (new_n9693_),
	   .A2 (new_n7276_),
	   .A1 (new_n7733_) );
   CLKBUF_X1 g2962 (
	   .Z (n4343),
	   .A (_net_7791) );
   CLKBUF_X1 g2961 (
	   .Z (n4338),
	   .A (_net_7808) );
   AND2_X1 g2960 (
	   .ZN (n4333),
	   .A2 (net_379),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g2959 (
	   .Z (n4330),
	   .A (net_6978) );
   CLKBUF_X1 g2958 (
	   .Z (n4326),
	   .A (net_6387) );
   NOR4_X1 g2957 (
	   .ZN (n4322),
	   .A4 (new_n8185_),
	   .A3 (new_n9686_),
	   .A2 (new_n9685_),
	   .A1 (new_n9684_) );
   NAND2_X1 g2956 (
	   .ZN (new_n9686_),
	   .A2 (_net_6404),
	   .A1 (new_n8186_) );
   INV_X1 g2955 (
	   .ZN (new_n9685_),
	   .A (new_n8265_) );
   NAND3_X1 g2954 (
	   .ZN (new_n9684_),
	   .A3 (new_n9304_),
	   .A2 (new_n9683_1_),
	   .A1 (new_n9682_) );
   INV_X1 g2953 (
	   .ZN (new_n9683_1_),
	   .A (_net_6405) );
   INV_X1 g2952 (
	   .ZN (new_n9682_),
	   .A (_net_6406) );
   CLKBUF_X1 g2951 (
	   .Z (n4318),
	   .A (net_6471) );
   OAI21_X1 g2950 (
	   .ZN (n4313),
	   .B2 (new_n9679_),
	   .B1 (new_n9674_),
	   .A (new_n9677_) );
   OAI21_X1 g2949 (
	   .ZN (new_n9679_),
	   .B2 (new_n9678_1_),
	   .B1 (n7691),
	   .A (new_n9440_) );
   NAND2_X1 g2948 (
	   .ZN (new_n9678_1_),
	   .A2 (_net_6422),
	   .A1 (new_n9676_) );
   NAND3_X1 g2947 (
	   .ZN (new_n9677_),
	   .A3 (new_n9676_),
	   .A2 (new_n9674_),
	   .A1 (new_n9673_1_) );
   NOR2_X1 g2946 (
	   .ZN (new_n9676_),
	   .A2 (new_n9435_),
	   .A1 (new_n9675_) );
   NAND3_X1 g2945 (
	   .ZN (new_n9675_),
	   .A3 (_net_6418),
	   .A2 (_net_6420),
	   .A1 (_net_6419) );
   INV_X1 g2944 (
	   .ZN (new_n9674_),
	   .A (_net_6422) );
   NOR2_X1 g2943 (
	   .ZN (new_n9673_1_),
	   .A2 (_net_6401),
	   .A1 (n7691) );
   CLKBUF_X1 g2942 (
	   .Z (n4309),
	   .A (net_6753) );
   NAND4_X1 g2941 (
	   .ZN (n4299),
	   .A4 (new_n9670_),
	   .A3 (new_n9666_),
	   .A2 (new_n9665_),
	   .A1 (new_n9664_1_) );
   NAND2_X1 g2940 (
	   .ZN (new_n9670_),
	   .A2 (new_n6879_),
	   .A1 (new_n9669_) );
   NAND2_X1 g2939 (
	   .ZN (new_n9669_),
	   .A2 (new_n9668_1_),
	   .A1 (new_n9667_) );
   AOI22_X1 g2938 (
	   .ZN (new_n9668_1_),
	   .B2 (net_6829),
	   .B1 (new_n6836_1_),
	   .A2 (net_6861),
	   .A1 (new_n6832_) );
   AOI22_X1 g2937 (
	   .ZN (new_n9667_),
	   .B2 (net_6925),
	   .B1 (new_n6873_),
	   .A2 (new_n6840_1_),
	   .A1 (net_6893) );
   NAND2_X1 g2936 (
	   .ZN (new_n9666_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n9249_) );
   NAND2_X1 g2935 (
	   .ZN (new_n9665_),
	   .A2 (new_n9178_1_),
	   .A1 (new_n9255_) );
   AOI22_X1 g2934 (
	   .ZN (new_n9664_1_),
	   .B2 (new_n6869_),
	   .B1 (_net_6128),
	   .A2 (new_n6854_),
	   .A1 (new_n9253_) );
   OAI21_X1 g2933 (
	   .ZN (n4294),
	   .B2 (new_n7225_),
	   .B1 (new_n9662_),
	   .A (new_n9661_) );
   INV_X1 g2932 (
	   .ZN (new_n9662_),
	   .A (_net_7318) );
   NAND2_X1 g2931 (
	   .ZN (new_n9661_),
	   .A2 (new_n9002_),
	   .A1 (new_n7222_) );
   XNOR2_X1 g2930 (
	   .ZN (n4289),
	   .B (new_n9659_),
	   .A (new_n8957_) );
   NAND2_X1 g2929 (
	   .ZN (new_n9659_),
	   .A2 (net_7529),
	   .A1 (new_n7268_) );
   CLKBUF_X1 g2928 (
	   .Z (n4284),
	   .A (x1459) );
   CLKBUF_X1 g2927 (
	   .Z (n4280),
	   .A (_net_7794) );
   CLKBUF_X1 g2926 (
	   .Z (n4271),
	   .A (net_6387) );
   CLKBUF_X1 g2925 (
	   .Z (n4267),
	   .A (_net_7796) );
   CLKBUF_X1 g2924 (
	   .Z (n4258),
	   .A (_net_7816) );
   CLKBUF_X1 g2923 (
	   .Z (n4253),
	   .A (net_6391) );
   NAND3_X1 g2922 (
	   .ZN (n4249),
	   .A3 (new_n9651_1_),
	   .A2 (new_n9650_),
	   .A1 (new_n9646_) );
   AOI22_X1 g2921 (
	   .ZN (new_n9651_1_),
	   .B2 (new_n8180_),
	   .B1 (net_7080),
	   .A2 (new_n7060_),
	   .A1 (new_n7065_) );
   AND3_X1 g2920 (
	   .ZN (new_n9650_),
	   .A3 (new_n9649_),
	   .A2 (new_n9648_),
	   .A1 (new_n9647_1_) );
   NAND2_X1 g2919 (
	   .ZN (new_n9649_),
	   .A2 (_net_6152),
	   .A1 (new_n7092_) );
   NAND2_X1 g2918 (
	   .ZN (new_n9648_),
	   .A2 (new_n7070_),
	   .A1 (new_n7086_) );
   NAND2_X1 g2917 (
	   .ZN (new_n9647_1_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n8845_1_) );
   AND3_X1 g2916 (
	   .ZN (new_n9646_),
	   .A3 (new_n9645_),
	   .A2 (new_n9644_),
	   .A1 (new_n9643_) );
   NAND4_X1 g2915 (
	   .ZN (new_n9645_),
	   .A4 (new_n7044_),
	   .A3 (_net_7092),
	   .A2 (net_7048),
	   .A1 (new_n8158_) );
   NAND4_X1 g2914 (
	   .ZN (new_n9644_),
	   .A4 (new_n7052_),
	   .A3 (net_6984),
	   .A2 (_net_7092),
	   .A1 (new_n8158_) );
   NAND4_X1 g2913 (
	   .ZN (new_n9643_),
	   .A4 (new_n7050_),
	   .A3 (_net_7092),
	   .A2 (net_7016),
	   .A1 (new_n8155_) );
   CLKBUF_X1 g2912 (
	   .Z (n4245),
	   .A (net_7398) );
   MUX2_X1 g2911 (
	   .Z (n4240),
	   .S (new_n7504_),
	   .B (_net_7635),
	   .A (new_n7216_1_) );
   CLKBUF_X1 g2910 (
	   .Z (n4235),
	   .A (_net_7813) );
   CLKBUF_X1 g2909 (
	   .Z (n4231),
	   .A (net_5858) );
   NOR2_X1 g2908 (
	   .ZN (n4226),
	   .A2 (new_n9637_),
	   .A1 (new_n9630_) );
   NAND4_X1 g2907 (
	   .ZN (new_n9637_),
	   .A4 (new_n9636_),
	   .A3 (new_n9634_),
	   .A2 (new_n9633_1_),
	   .A1 (new_n9631_) );
   NAND2_X1 g2906 (
	   .ZN (new_n9636_),
	   .A2 (_net_6827),
	   .A1 (new_n9635_) );
   NAND2_X1 g2905 (
	   .ZN (new_n9635_),
	   .A2 (new_n9627_),
	   .A1 (new_n9632_) );
   OAI21_X1 g2904 (
	   .ZN (new_n9634_),
	   .B2 (new_n8389_),
	   .B1 (new_n8394_),
	   .A (new_n7554_) );
   NAND3_X1 g2903 (
	   .ZN (new_n9633_1_),
	   .A3 (new_n9627_),
	   .A2 (new_n8303_1_),
	   .A1 (new_n9632_) );
   OAI21_X1 g2902 (
	   .ZN (new_n9632_),
	   .B2 (new_n7570_),
	   .B1 (new_n7554_),
	   .A (new_n7568_) );
   OAI21_X1 g2901 (
	   .ZN (new_n9631_),
	   .B2 (new_n8764_),
	   .B1 (n2948),
	   .A (_net_6822) );
   XNOR2_X1 g2900 (
	   .ZN (new_n9630_),
	   .B (new_n9629_),
	   .A (new_n9628_1_) );
   INV_X1 g2899 (
	   .ZN (new_n9629_),
	   .A (_net_6828) );
   XNOR2_X1 g2898 (
	   .ZN (new_n9628_1_),
	   .B (_net_6825),
	   .A (new_n9627_) );
   NAND3_X1 g2897 (
	   .ZN (new_n9627_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (_net_6822) );
   CLKBUF_X1 g2896 (
	   .Z (n4221),
	   .A (_net_7814) );
   MUX2_X1 g2895 (
	   .Z (n4217),
	   .S (new_n7504_),
	   .B (_net_7630),
	   .A (new_n9405_1_) );
   OAI221_X1 g2894 (
	   .ZN (n4212),
	   .C2 (new_n7306_),
	   .C1 (new_n9517_1_),
	   .B2 (new_n7303_),
	   .B1 (new_n9039_),
	   .A (new_n9623_) );
   AOI22_X1 g2893 (
	   .ZN (new_n9623_),
	   .B2 (_net_7414),
	   .B1 (new_n9203_),
	   .A2 (_net_7446),
	   .A1 (new_n8694_1_) );
   CLKBUF_X1 g2892 (
	   .Z (n4207),
	   .A (_net_7808) );
   OAI21_X1 g2891 (
	   .ZN (n4203),
	   .B2 (new_n9620_1_),
	   .B1 (new_n9619_),
	   .A (new_n9618_) );
   INV_X1 g2890 (
	   .ZN (new_n9620_1_),
	   .A (_net_189) );
   INV_X1 g2889 (
	   .ZN (new_n9619_),
	   .A (new_n6941_) );
   INV_X1 g2888 (
	   .ZN (new_n9618_),
	   .A (_net_277) );
   CLKBUF_X1 g2887 (
	   .Z (n4199),
	   .A (net_6447) );
   CLKBUF_X1 g2886 (
	   .Z (n4194),
	   .A (_net_7822) );
   CLKBUF_X1 g2885 (
	   .Z (n4191),
	   .A (net_7123) );
   OAI21_X1 g2884 (
	   .ZN (n4186),
	   .B2 (new_n7225_),
	   .B1 (new_n9613_),
	   .A (new_n9612_) );
   INV_X1 g2883 (
	   .ZN (new_n9613_),
	   .A (_net_7321) );
   NAND2_X1 g2882 (
	   .ZN (new_n9612_),
	   .A2 (new_n9611_1_),
	   .A1 (new_n7222_) );
   OAI221_X1 g2881 (
	   .ZN (new_n9611_1_),
	   .C2 (new_n7107_1_),
	   .C1 (new_n7105_),
	   .B2 (new_n8132_),
	   .B1 (new_n7106_),
	   .A (new_n9610_) );
   NAND2_X1 g2880 (
	   .ZN (new_n9610_),
	   .A2 (net_7241),
	   .A1 (new_n6942_) );
   NAND2_X1 g2879 (
	   .ZN (n4181),
	   .A2 (new_n9608_),
	   .A1 (new_n9607_) );
   AOI22_X1 g2878 (
	   .ZN (new_n9608_),
	   .B2 (_net_7556),
	   .B1 (new_n6755_),
	   .A2 (_net_7620),
	   .A1 (new_n6746_1_) );
   AOI22_X1 g2877 (
	   .ZN (new_n9607_),
	   .B2 (_net_7588),
	   .B1 (new_n7350_),
	   .A2 (new_n7970_1_),
	   .A1 (_net_7652) );
   CLKBUF_X1 g2876 (
	   .Z (n4176),
	   .A (_net_6087) );
   INV_X1 g2875 (
	   .ZN (n4171),
	   .A (new_n9604_) );
   NAND2_X1 g2874 (
	   .ZN (new_n9604_),
	   .A2 (new_n9420_1_),
	   .A1 (new_n7448_) );
   OAI21_X1 g2873 (
	   .ZN (n4166),
	   .B2 (new_n7279_),
	   .B1 (new_n9602_1_),
	   .A (new_n9601_) );
   INV_X1 g2872 (
	   .ZN (new_n9602_1_),
	   .A (_net_7437) );
   NAND2_X1 g2871 (
	   .ZN (new_n9601_),
	   .A2 (new_n8859_),
	   .A1 (new_n7272_) );
   CLKBUF_X1 g2870 (
	   .Z (n4161),
	   .A (net_6382) );
   CLKBUF_X1 g2869 (
	   .Z (n4158),
	   .A (net_6714) );
   CLKBUF_X1 g2868 (
	   .Z (n4153),
	   .A (net_145) );
   CLKBUF_X1 g2867 (
	   .Z (n4148),
	   .A (_net_7793) );
   CLKBUF_X1 g2866 (
	   .Z (n4145),
	   .A (net_6592) );
   OAI21_X1 g2865 (
	   .ZN (n4140),
	   .B2 (new_n7111_1_),
	   .B1 (new_n9594_),
	   .A (new_n9593_) );
   INV_X1 g2864 (
	   .ZN (new_n9594_),
	   .A (_net_7347) );
   NAND2_X1 g2863 (
	   .ZN (new_n9593_),
	   .A2 (new_n7773_1_),
	   .A1 (new_n7101_) );
   NOR3_X1 g2862 (
	   .ZN (n4135),
	   .A3 (new_n8754_),
	   .A2 (new_n9591_),
	   .A1 (new_n9590_) );
   AOI21_X1 g2861 (
	   .ZN (new_n9591_),
	   .B2 (_net_5983),
	   .B1 (net_7231),
	   .A (_net_7232) );
   AND3_X1 g2860 (
	   .ZN (new_n9590_),
	   .A3 (_net_5983),
	   .A2 (_net_7232),
	   .A1 (net_7231) );
   CLKBUF_X1 g2859 (
	   .Z (n4131),
	   .A (net_7400) );
   AOI21_X1 g2858 (
	   .ZN (n4126),
	   .B2 (new_n9586_),
	   .B1 (new_n8025_),
	   .A (new_n9587_) );
   OAI21_X1 g2857 (
	   .ZN (new_n9587_),
	   .B2 (new_n8025_),
	   .B1 (new_n9586_),
	   .A (_net_6039) );
   NAND3_X1 g2856 (
	   .ZN (new_n9586_),
	   .A3 (new_n7810_1_),
	   .A2 (new_n7686_1_),
	   .A1 (n1600) );
   OAI21_X1 g2855 (
	   .ZN (n4121),
	   .B2 (new_n9351_),
	   .B1 (new_n9584_),
	   .A (new_n9583_1_) );
   INV_X1 g2854 (
	   .ZN (new_n9584_),
	   .A (_net_188) );
   INV_X1 g2853 (
	   .ZN (new_n9583_1_),
	   .A (_net_276) );
   OAI21_X1 g2852 (
	   .ZN (n4116),
	   .B2 (new_n7111_1_),
	   .B1 (new_n9581_),
	   .A (new_n9580_) );
   INV_X1 g2851 (
	   .ZN (new_n9581_),
	   .A (_net_7364) );
   NAND2_X1 g2850 (
	   .ZN (new_n9580_),
	   .A2 (new_n7335_1_),
	   .A1 (new_n7101_) );
   CLKBUF_X1 g2849 (
	   .Z (n4112),
	   .A (net_6867) );
   MUX2_X1 g2848 (
	   .Z (n4107),
	   .S (new_n7285_),
	   .B (_net_7719),
	   .A (_net_7821) );
   CLKBUF_X1 g2847 (
	   .Z (n4102),
	   .A (_net_7813) );
   CLKBUF_X1 g2846 (
	   .Z (n4098),
	   .A (_net_7798) );
   OAI21_X1 g2845 (
	   .ZN (n4094),
	   .B2 (new_n7652_),
	   .B1 (new_n9574_1_),
	   .A (new_n9573_) );
   INV_X1 g2844 (
	   .ZN (new_n9574_1_),
	   .A (_net_7404) );
   NAND2_X1 g2843 (
	   .ZN (new_n9573_),
	   .A2 (new_n8066_),
	   .A1 (new_n7646_) );
   NAND3_X1 g2842 (
	   .ZN (n4089),
	   .A3 (new_n9571_),
	   .A2 (new_n6963_),
	   .A1 (new_n9570_) );
   NAND2_X1 g2841 (
	   .ZN (new_n9571_),
	   .A2 (new_n8183_1_),
	   .A1 (new_n9569_1_) );
   OR2_X1 g2840 (
	   .ZN (new_n9570_),
	   .A2 (new_n8183_1_),
	   .A1 (new_n9569_1_) );
   AND4_X1 g2839 (
	   .ZN (new_n9569_1_),
	   .A4 (_net_6409),
	   .A3 (_net_6410),
	   .A2 (new_n9305_),
	   .A1 (_net_6408) );
   MUX2_X1 g2838 (
	   .Z (n4084),
	   .S (new_n7538_),
	   .B (_net_294),
	   .A (_net_7814) );
   AND2_X1 g2837 (
	   .ZN (n4079),
	   .A2 (net_374),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g2836 (
	   .Z (n4075),
	   .A (net_6399) );
   CLKBUF_X1 g2835 (
	   .Z (n4071),
	   .A (_net_7814) );
   CLKBUF_X1 g2834 (
	   .Z (n4068),
	   .A (net_6444) );
   OAI21_X1 g2833 (
	   .ZN (n4063),
	   .B2 (new_n7225_),
	   .B1 (new_n9562_),
	   .A (new_n9561_) );
   INV_X1 g2832 (
	   .ZN (new_n9562_),
	   .A (_net_7329) );
   NAND2_X1 g2831 (
	   .ZN (new_n9561_),
	   .A2 (new_n9560_),
	   .A1 (new_n7222_) );
   OAI21_X1 g2830 (
	   .ZN (new_n9560_),
	   .B2 (new_n9559_1_),
	   .B1 (new_n6951_),
	   .A (new_n9558_) );
   INV_X1 g2829 (
	   .ZN (new_n9559_1_),
	   .A (net_7249) );
   AOI22_X1 g2828 (
	   .ZN (new_n9558_),
	   .B2 (_net_269),
	   .B1 (net_343),
	   .A2 (net_341),
	   .A1 (_net_270) );
   CLKBUF_X1 g2827 (
	   .Z (n4059),
	   .A (net_7013) );
   CLKBUF_X1 g2826 (
	   .Z (n4055),
	   .A (net_7711) );
   CLKBUF_X1 g2825 (
	   .Z (n4051),
	   .A (net_6613) );
   CLKBUF_X1 g2824 (
	   .Z (n4046),
	   .A (net_6390) );
   MUX2_X1 g2823 (
	   .Z (n4042),
	   .S (new_n7504_),
	   .B (_net_7633),
	   .A (new_n9349_) );
   CLKBUF_X1 g2822 (
	   .Z (n4037),
	   .A (_net_7793) );
   CLKBUF_X1 g2821 (
	   .Z (n4033),
	   .A (_net_7821) );
   MUX2_X1 g2820 (
	   .Z (n4029),
	   .S (new_n7029_),
	   .B (_net_7601),
	   .A (new_n9349_) );
   CLKBUF_X1 g2819 (
	   .Z (n4024),
	   .A (_net_7804) );
   CLKBUF_X1 g2818 (
	   .Z (n4020),
	   .A (_net_7813) );
   AOI21_X1 g2817 (
	   .ZN (n4016),
	   .B2 (new_n9546_1_),
	   .B1 (new_n8424_),
	   .A (new_n7428_) );
   INV_X1 g2816 (
	   .ZN (new_n9546_1_),
	   .A (_net_6027) );
   CLKBUF_X1 g2815 (
	   .Z (n4011),
	   .A (_net_6103) );
   CLKBUF_X1 g2814 (
	   .Z (n4007),
	   .A (net_6852) );
   CLKBUF_X1 g2813 (
	   .Z (n4002),
	   .A (_net_7817) );
   NAND2_X1 g2812 (
	   .ZN (n3998),
	   .A2 (new_n9541_1_),
	   .A1 (new_n9538_) );
   NAND3_X1 g2811 (
	   .ZN (new_n9541_1_),
	   .A3 (new_n9540_),
	   .A2 (new_n9539_),
	   .A1 (new_n7287_) );
   NAND2_X1 g2810 (
	   .ZN (new_n9540_),
	   .A2 (new_n8921_),
	   .A1 (new_n7045_1_) );
   INV_X1 g2809 (
	   .ZN (new_n9539_),
	   .A (new_n9536_) );
   AOI22_X1 g2808 (
	   .ZN (new_n9538_),
	   .B2 (_net_7095),
	   .B1 (new_n7092_),
	   .A2 (new_n8155_),
	   .A1 (new_n9537_1_) );
   AOI22_X1 g2807 (
	   .ZN (new_n9537_1_),
	   .B2 (new_n7290_),
	   .B1 (new_n8921_),
	   .A2 (_net_7092),
	   .A1 (new_n9536_) );
   NOR2_X1 g2806 (
	   .ZN (new_n9536_),
	   .A2 (new_n8921_),
	   .A1 (new_n7045_1_) );
   CLKBUF_X1 g2805 (
	   .Z (n3993),
	   .A (_net_7795) );
   CLKBUF_X1 g2804 (
	   .Z (n3989),
	   .A (net_6392) );
   CLKBUF_X1 g2803 (
	   .Z (n3985),
	   .A (_net_7815) );
   NAND2_X1 g2802 (
	   .ZN (n3981),
	   .A2 (new_n9531_),
	   .A1 (new_n9526_) );
   AND4_X1 g2801 (
	   .ZN (new_n9531_),
	   .A4 (new_n9530_),
	   .A3 (new_n9529_),
	   .A2 (new_n9528_1_),
	   .A1 (new_n9527_) );
   NAND2_X1 g2800 (
	   .ZN (new_n9530_),
	   .A2 (_net_6112),
	   .A1 (new_n7210_) );
   NAND2_X1 g2799 (
	   .ZN (new_n9529_),
	   .A2 (new_n7587_),
	   .A1 (new_n9032_) );
   NAND2_X1 g2798 (
	   .ZN (new_n9528_1_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n9493_) );
   NAND2_X1 g2797 (
	   .ZN (new_n9527_),
	   .A2 (new_n8252_),
	   .A1 (new_n7565_) );
   AND4_X1 g2796 (
	   .ZN (new_n9526_),
	   .A4 (new_n9525_1_),
	   .A3 (new_n9524_),
	   .A2 (new_n9523_),
	   .A1 (new_n9522_) );
   NAND4_X1 g2795 (
	   .ZN (new_n9525_1_),
	   .A4 (new_n7194_1_),
	   .A3 (_net_6822),
	   .A2 (net_6746),
	   .A1 (new_n7559_) );
   NAND4_X1 g2794 (
	   .ZN (new_n9524_),
	   .A4 (new_n7191_),
	   .A3 (net_6778),
	   .A2 (_net_6822),
	   .A1 (new_n7560_) );
   NAND3_X1 g2793 (
	   .ZN (new_n9523_),
	   .A3 (new_n7189_),
	   .A2 (net_6810),
	   .A1 (new_n7555_) );
   NAND3_X1 g2792 (
	   .ZN (new_n9522_),
	   .A3 (new_n7196_),
	   .A2 (net_6714),
	   .A1 (new_n7556_) );
   AND2_X1 g2791 (
	   .ZN (n3976),
	   .A2 (_net_6201),
	   .A1 (new_n9520_1_) );
   BUF_X2 g2790 (
	   .Z (new_n9520_1_),
	   .A (new_n7235_1_) );
   CLKBUF_X1 g2789 (
	   .Z (n3972),
	   .A (net_7537) );
   OAI21_X1 g2788 (
	   .ZN (n3967),
	   .B2 (new_n7736_),
	   .B1 (new_n9517_1_),
	   .A (new_n9516_) );
   INV_X1 g2787 (
	   .ZN (new_n9517_1_),
	   .A (_net_7510) );
   NAND2_X1 g2786 (
	   .ZN (new_n9516_),
	   .A2 (new_n9037_1_),
	   .A1 (new_n7733_) );
   CLKBUF_X1 g2785 (
	   .Z (n3962),
	   .A (_net_6176) );
   CLKBUF_X1 g2784 (
	   .Z (n3957),
	   .A (net_6387) );
   CLKBUF_X1 g2783 (
	   .Z (n3953),
	   .A (_net_7815) );
   CLKBUF_X1 g2782 (
	   .Z (n3949),
	   .A (_net_7822) );
   CLKBUF_X1 g2781 (
	   .Z (n3945),
	   .A (net_6384) );
   MUX2_X1 g2780 (
	   .Z (n3941),
	   .S (new_n7029_),
	   .B (_net_7591),
	   .A (new_n9509_) );
   OAI21_X1 g2779 (
	   .ZN (new_n9509_),
	   .B2 (new_n9508_),
	   .B1 (new_n7019_),
	   .A (new_n9507_1_) );
   INV_X1 g2778 (
	   .ZN (new_n9508_),
	   .A (net_7543) );
   AOI22_X1 g2777 (
	   .ZN (new_n9507_1_),
	   .B2 (_net_291),
	   .B1 (net_375),
	   .A2 (_net_292),
	   .A1 (net_373) );
   CLKBUF_X1 g2776 (
	   .Z (n3936),
	   .A (_net_7823) );
   OAI21_X1 g2775 (
	   .ZN (n3932),
	   .B2 (new_n7652_),
	   .B1 (new_n9504_),
	   .A (new_n9503_) );
   INV_X1 g2774 (
	   .ZN (new_n9504_),
	   .A (_net_7418) );
   NAND2_X1 g2773 (
	   .ZN (new_n9503_),
	   .A2 (new_n9502_1_),
	   .A1 (new_n7646_) );
   OAI21_X1 g2772 (
	   .ZN (new_n9502_1_),
	   .B2 (new_n7961_),
	   .B1 (new_n7034_),
	   .A (new_n9501_) );
   AOI22_X1 g2771 (
	   .ZN (new_n9501_),
	   .B2 (_net_281),
	   .B1 (net_363),
	   .A2 (_net_280),
	   .A1 (net_365) );
   MUX2_X1 g2770 (
	   .Z (n3927),
	   .S (new_n7609_),
	   .B (_net_7563),
	   .A (new_n7022_) );
   NAND2_X1 g2769 (
	   .ZN (n3922),
	   .A2 (new_n9498_),
	   .A1 (new_n9488_) );
   AND4_X1 g2768 (
	   .ZN (new_n9498_),
	   .A4 (new_n9497_1_),
	   .A3 (new_n9496_),
	   .A2 (new_n9495_),
	   .A1 (new_n9494_) );
   NAND2_X1 g2767 (
	   .ZN (new_n9497_1_),
	   .A2 (_net_6116),
	   .A1 (new_n7210_) );
   NAND2_X1 g2766 (
	   .ZN (new_n9496_),
	   .A2 (new_n7587_),
	   .A1 (new_n8617_) );
   NAND2_X1 g2765 (
	   .ZN (new_n9495_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n7573_) );
   NAND2_X1 g2764 (
	   .ZN (new_n9494_),
	   .A2 (new_n9493_),
	   .A1 (new_n7565_) );
   NAND4_X1 g2763 (
	   .ZN (new_n9493_),
	   .A4 (new_n9492_1_),
	   .A3 (new_n9491_),
	   .A2 (new_n9490_),
	   .A1 (new_n9489_) );
   NAND3_X1 g2762 (
	   .ZN (new_n9492_1_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6798) );
   NAND3_X1 g2761 (
	   .ZN (new_n9491_),
	   .A3 (_net_6824),
	   .A2 (net_6766),
	   .A1 (new_n7570_) );
   NAND3_X1 g2760 (
	   .ZN (new_n9490_),
	   .A3 (_net_6823),
	   .A2 (net_6734),
	   .A1 (new_n7568_) );
   NAND2_X1 g2759 (
	   .ZN (new_n9489_),
	   .A2 (net_6702),
	   .A1 (new_n7566_) );
   AND4_X1 g2758 (
	   .ZN (new_n9488_),
	   .A4 (new_n9487_1_),
	   .A3 (new_n9486_),
	   .A2 (new_n9485_),
	   .A1 (new_n9484_) );
   NAND4_X1 g2757 (
	   .ZN (new_n9487_1_),
	   .A4 (new_n7194_1_),
	   .A3 (net_6750),
	   .A2 (_net_6822),
	   .A1 (new_n7559_) );
   NAND4_X1 g2756 (
	   .ZN (new_n9486_),
	   .A4 (new_n7191_),
	   .A3 (net_6782),
	   .A2 (_net_6822),
	   .A1 (new_n7560_) );
   NAND3_X1 g2755 (
	   .ZN (new_n9485_),
	   .A3 (new_n7189_),
	   .A2 (net_6814),
	   .A1 (new_n7555_) );
   NAND3_X1 g2754 (
	   .ZN (new_n9484_),
	   .A3 (new_n7196_),
	   .A2 (net_6718),
	   .A1 (new_n7556_) );
   CLKBUF_X1 g2753 (
	   .Z (n3917),
	   .A (_net_7814) );
   AOI21_X1 g2752 (
	   .ZN (n3913),
	   .B2 (new_n7326_1_),
	   .B1 (new_n9481_),
	   .A (new_n9480_) );
   INV_X1 g2751 (
	   .ZN (new_n9481_),
	   .A (_net_7270) );
   NOR2_X1 g2750 (
	   .ZN (new_n9480_),
	   .A2 (n1029),
	   .A1 (new_n7325_) );
   NAND2_X1 g2749 (
	   .ZN (n3908),
	   .A2 (new_n9478_1_),
	   .A1 (new_n9477_) );
   AOI22_X1 g2748 (
	   .ZN (new_n9478_1_),
	   .B2 (net_7527),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7495) );
   AOI22_X1 g2747 (
	   .ZN (new_n9477_),
	   .B2 (_net_7431),
	   .B1 (new_n7298_),
	   .A2 (net_7463),
	   .A1 (new_n7296_) );
   CLKBUF_X1 g2746 (
	   .Z (n3904),
	   .A (net_7239) );
   CLKBUF_X1 g2745 (
	   .Z (n3899),
	   .A (net_7799) );
   CLKBUF_X1 g2744 (
	   .Z (n3896),
	   .A (net_6855) );
   MUX2_X1 g2743 (
	   .Z (n3891),
	   .S (_net_154),
	   .B (net_319),
	   .A (_net_123) );
   MUX2_X1 g2742 (
	   .Z (n3886),
	   .S (new_n7609_),
	   .B (_net_7574),
	   .A (n2850) );
   CLKBUF_X1 g2741 (
	   .Z (n3881),
	   .A (net_7799) );
   OAI21_X1 g2740 (
	   .ZN (n3877),
	   .B2 (new_n9469_),
	   .B1 (new_n9468_),
	   .A (new_n9467_1_) );
   INV_X1 g2739 (
	   .ZN (new_n9469_),
	   .A (new_n6813_1_) );
   INV_X1 g2738 (
	   .ZN (new_n9468_),
	   .A (_net_6065) );
   NAND2_X1 g2737 (
	   .ZN (new_n9467_1_),
	   .A2 (new_n7166_),
	   .A1 (new_n8146_) );
   NOR3_X1 g2736 (
	   .ZN (n3872),
	   .A3 (new_n6944_),
	   .A2 (new_n9465_),
	   .A1 (new_n9463_) );
   INV_X1 g2735 (
	   .ZN (new_n9465_),
	   .A (new_n9464_) );
   XNOR2_X1 g2734 (
	   .ZN (new_n9464_),
	   .B (_net_7384),
	   .A (_net_7380) );
   NAND2_X1 g2733 (
	   .ZN (new_n9463_),
	   .A2 (new_n9462_1_),
	   .A1 (n3464) );
   XNOR2_X1 g2732 (
	   .ZN (new_n9462_1_),
	   .B (_net_7383),
	   .A (_net_7379) );
   CLKBUF_X1 g2731 (
	   .Z (n3867),
	   .A (_net_7806) );
   CLKBUF_X1 g2730 (
	   .Z (n3864),
	   .A (net_6850) );
   OAI21_X1 g2729 (
	   .ZN (n3859),
	   .B2 (new_n7258_),
	   .B1 (new_n9458_),
	   .A (new_n9457_) );
   INV_X1 g2728 (
	   .ZN (new_n9458_),
	   .A (_net_7290) );
   NAND2_X1 g2727 (
	   .ZN (new_n9457_),
	   .A2 (new_n7495_),
	   .A1 (new_n7252_1_) );
   CLKBUF_X1 g2726 (
	   .Z (n3855),
	   .A (net_6595) );
   CLKBUF_X1 g2725 (
	   .Z (n3851),
	   .A (net_6829) );
   NAND3_X1 g2724 (
	   .ZN (n3846),
	   .A3 (new_n9453_),
	   .A2 (new_n9452_),
	   .A1 (new_n9448_) );
   AOI22_X1 g2723 (
	   .ZN (new_n9453_),
	   .B2 (new_n8180_),
	   .B1 (net_7086),
	   .A2 (new_n8837_),
	   .A1 (new_n7060_) );
   AND3_X1 g2722 (
	   .ZN (new_n9452_),
	   .A3 (new_n9451_),
	   .A2 (new_n9450_),
	   .A1 (new_n9449_1_) );
   NAND2_X1 g2721 (
	   .ZN (new_n9451_),
	   .A2 (_net_6158),
	   .A1 (new_n7092_) );
   NAND2_X1 g2720 (
	   .ZN (new_n9450_),
	   .A2 (new_n7070_),
	   .A1 (new_n8670_) );
   NAND2_X1 g2719 (
	   .ZN (new_n9449_1_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n8662_1_) );
   AND3_X1 g2718 (
	   .ZN (new_n9448_),
	   .A3 (new_n9447_),
	   .A2 (new_n9446_),
	   .A1 (new_n9445_1_) );
   NAND4_X1 g2717 (
	   .ZN (new_n9447_),
	   .A4 (new_n7044_),
	   .A3 (net_7054),
	   .A2 (_net_7092),
	   .A1 (new_n8158_) );
   NAND4_X1 g2716 (
	   .ZN (new_n9446_),
	   .A4 (new_n7052_),
	   .A3 (net_6990),
	   .A2 (_net_7092),
	   .A1 (new_n8158_) );
   NAND4_X1 g2715 (
	   .ZN (new_n9445_1_),
	   .A4 (new_n7050_),
	   .A3 (_net_7092),
	   .A2 (net_7022),
	   .A1 (new_n8155_) );
   MUX2_X1 g2714 (
	   .Z (n3841),
	   .S (new_n7545_),
	   .B (_net_7652),
	   .A (new_n8475_) );
   AOI21_X1 g2713 (
	   .ZN (n3836),
	   .B2 (new_n9442_),
	   .B1 (_net_6419),
	   .A (new_n9441_1_) );
   NOR2_X1 g2712 (
	   .ZN (new_n9442_),
	   .A2 (new_n9438_),
	   .A1 (n7691) );
   NAND2_X1 g2711 (
	   .ZN (new_n9441_1_),
	   .A2 (new_n9440_),
	   .A1 (new_n9439_) );
   INV_X1 g2710 (
	   .ZN (new_n9440_),
	   .A (_net_6401) );
   OAI21_X1 g2709 (
	   .ZN (new_n9439_),
	   .B2 (new_n9438_),
	   .B1 (n7691),
	   .A (new_n9433_) );
   INV_X1 g2708 (
	   .ZN (new_n9438_),
	   .A (_net_6418) );
   NOR3_X1 g2707 (
	   .ZN (n7691),
	   .A3 (_net_6422),
	   .A2 (_net_6419),
	   .A1 (new_n9436_1_) );
   NAND4_X1 g2706 (
	   .ZN (new_n9436_1_),
	   .A4 (_net_6418),
	   .A3 (_net_6423),
	   .A2 (new_n9435_),
	   .A1 (new_n9434_) );
   INV_X1 g2705 (
	   .ZN (new_n9435_),
	   .A (_net_6421) );
   INV_X1 g2704 (
	   .ZN (new_n9434_),
	   .A (_net_6420) );
   INV_X1 g2703 (
	   .ZN (new_n9433_),
	   .A (_net_6419) );
   CLKBUF_X1 g2702 (
	   .Z (n3831),
	   .A (net_7802) );
   CLKBUF_X1 g2701 (
	   .Z (n3822),
	   .A (_net_6076) );
   CLKBUF_X1 g2700 (
	   .Z (n3817),
	   .A (net_6394) );
   OAI221_X1 g2699 (
	   .ZN (n3813),
	   .C2 (new_n6920_),
	   .C1 (new_n9428_1_),
	   .B2 (new_n6917_),
	   .B1 (new_n9427_),
	   .A (new_n9426_) );
   INV_X1 g2698 (
	   .ZN (new_n9428_1_),
	   .A (net_7372) );
   INV_X1 g2697 (
	   .ZN (new_n9427_),
	   .A (net_7308) );
   AOI22_X1 g2696 (
	   .ZN (new_n9426_),
	   .B2 (_net_7276),
	   .B1 (new_n6913_),
	   .A2 (net_7340),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g2695 (
	   .Z (n3809),
	   .A (net_6429) );
   CLKBUF_X1 g2694 (
	   .Z (n3805),
	   .A (net_7714) );
   CLKBUF_X1 g2693 (
	   .Z (n3801),
	   .A (net_7149) );
   AOI21_X1 g2692 (
	   .ZN (n3796),
	   .B2 (new_n9421_),
	   .B1 (new_n7446_1_),
	   .A (new_n7449_) );
   NAND2_X1 g2691 (
	   .ZN (new_n9421_),
	   .A2 (_net_7785),
	   .A1 (new_n9420_1_) );
   INV_X1 g2690 (
	   .ZN (new_n9420_1_),
	   .A (_net_7784) );
   CLKBUF_X1 g2689 (
	   .Z (n3791),
	   .A (_net_7804) );
   AOI21_X1 g2688 (
	   .ZN (n3787),
	   .B2 (new_n9416_),
	   .B1 (new_n7072_1_),
	   .A (new_n9417_) );
   OAI21_X1 g2687 (
	   .ZN (new_n9417_),
	   .B2 (new_n7072_1_),
	   .B1 (new_n9416_),
	   .A (_net_6028) );
   NAND2_X1 g2686 (
	   .ZN (new_n9416_),
	   .A2 (new_n7057_),
	   .A1 (new_n7056_) );
   MUX2_X1 g2685 (
	   .Z (n3782),
	   .S (new_n7504_),
	   .B (_net_7626),
	   .A (new_n7806_1_) );
   CLKBUF_X1 g2684 (
	   .Z (n3777),
	   .A (_net_7798) );
   CLKBUF_X1 g2683 (
	   .Z (n3773),
	   .A (_net_7796) );
   CLKBUF_X1 g2682 (
	   .Z (n3770),
	   .A (net_6991) );
   MUX2_X1 g2681 (
	   .Z (n3765),
	   .S (new_n7538_),
	   .B (_net_290),
	   .A (_net_7810) );
   CLKBUF_X1 g2680 (
	   .Z (n3761),
	   .A (net_6442) );
   CLKBUF_X1 g2679 (
	   .Z (n3756),
	   .A (net_6391) );
   CLKBUF_X1 g2678 (
	   .Z (n3752),
	   .A (_net_6069) );
   CLKBUF_X1 g2677 (
	   .Z (n3747),
	   .A (_net_6129) );
   MUX2_X1 g2676 (
	   .Z (n3742),
	   .S (new_n7029_),
	   .B (_net_7598),
	   .A (new_n9405_1_) );
   OAI21_X1 g2675 (
	   .ZN (new_n9405_1_),
	   .B2 (new_n9404_),
	   .B1 (new_n7019_),
	   .A (new_n9403_) );
   INV_X1 g2674 (
	   .ZN (new_n9404_),
	   .A (net_7550) );
   AOI22_X1 g2673 (
	   .ZN (new_n9403_),
	   .B2 (_net_291),
	   .B1 (net_382),
	   .A2 (_net_292),
	   .A1 (net_380) );
   OAI21_X1 g2672 (
	   .ZN (n3737),
	   .B2 (new_n7279_),
	   .B1 (new_n9401_),
	   .A (new_n9400_) );
   INV_X1 g2671 (
	   .ZN (new_n9401_),
	   .A (_net_7444) );
   NAND2_X1 g2670 (
	   .ZN (new_n9400_),
	   .A2 (new_n7649_1_),
	   .A1 (new_n7272_) );
   CLKBUF_X1 g2669 (
	   .Z (n3733),
	   .A (x1550) );
   CLKBUF_X1 g2668 (
	   .Z (n3729),
	   .A (_net_7813) );
   CLKBUF_X1 g2667 (
	   .Z (n3725),
	   .A (net_6881) );
   CLKBUF_X1 g2666 (
	   .Z (n3720),
	   .A (_net_6092) );
   CLKBUF_X1 g2665 (
	   .Z (n3716),
	   .A (net_6486) );
   AND2_X1 g2664 (
	   .ZN (n3711),
	   .A2 (new_n9393_1_),
	   .A1 (new_n9392_) );
   INV_X1 g2663 (
	   .ZN (new_n9393_1_),
	   .A (x977) );
   AOI211_X1 g2662 (
	   .ZN (new_n9392_),
	   .C2 (new_n7798_1_),
	   .C1 (new_n7797_),
	   .B (new_n6867_1_),
	   .A (new_n9391_) );
   INV_X1 g2661 (
	   .ZN (new_n9391_),
	   .A (_net_6023) );
   CLKBUF_X1 g2660 (
	   .Z (n3707),
	   .A (net_6721) );
   CLKBUF_X1 g2659 (
	   .Z (n3703),
	   .A (net_6976) );
   NOR2_X1 g2658 (
	   .ZN (n3698),
	   .A2 (x906),
	   .A1 (new_n9387_) );
   AOI21_X1 g2657 (
	   .ZN (new_n9387_),
	   .B2 (net_7777),
	   .B1 (new_n8760_),
	   .A (_net_5853) );
   OAI21_X1 g2656 (
	   .ZN (n3693),
	   .B2 (new_n6957_1_),
	   .B1 (new_n9385_1_),
	   .A (new_n9384_) );
   INV_X1 g2655 (
	   .ZN (new_n9385_1_),
	   .A (_net_7250) );
   NAND2_X1 g2654 (
	   .ZN (new_n9384_),
	   .A2 (new_n8780_1_),
	   .A1 (new_n6949_) );
   CLKBUF_X1 g2653 (
	   .Z (n3689),
	   .A (net_6605) );
   AOI21_X1 g2652 (
	   .ZN (n3684),
	   .B2 (new_n9381_1_),
	   .B1 (new_n9380_),
	   .A (x940) );
   INV_X1 g2651 (
	   .ZN (new_n9381_1_),
	   .A (_net_5854) );
   NAND3_X1 g2650 (
	   .ZN (new_n9380_),
	   .A3 (net_7776),
	   .A2 (_net_6034),
	   .A1 (n9592) );
   AOI21_X1 g2649 (
	   .ZN (n9592),
	   .B2 (new_n9378_),
	   .B1 (new_n9377_1_),
	   .A (new_n7090_) );
   AOI21_X1 g2648 (
	   .ZN (new_n9378_),
	   .B2 (new_n9376_),
	   .B1 (new_n9375_),
	   .A (_net_5976) );
   OAI21_X1 g2647 (
	   .ZN (new_n9377_1_),
	   .B2 (new_n9376_),
	   .B1 (new_n9375_),
	   .A (new_n9374_) );
   INV_X1 g2646 (
	   .ZN (new_n9376_),
	   .A (_net_5978) );
   NOR2_X1 g2645 (
	   .ZN (new_n9375_),
	   .A2 (_net_5977),
	   .A1 (_net_6032) );
   INV_X1 g2644 (
	   .ZN (new_n9374_),
	   .A (_net_6033) );
   CLKBUF_X1 g2643 (
	   .Z (n3679),
	   .A (_net_7801) );
   AOI21_X1 g2642 (
	   .ZN (n3675),
	   .B2 (new_n9371_),
	   .B1 (new_n9370_1_),
	   .A (new_n7428_) );
   INV_X1 g2641 (
	   .ZN (new_n9371_),
	   .A (_net_7728) );
   INV_X1 g2640 (
	   .ZN (new_n9370_1_),
	   .A (net_6014) );
   CLKBUF_X1 g2639 (
	   .Z (n3670),
	   .A (_net_7794) );
   AOI21_X1 g2638 (
	   .ZN (n3666),
	   .B2 (new_n7739_),
	   .B1 (new_n9367_),
	   .A (new_n9366_) );
   INV_X1 g2637 (
	   .ZN (new_n9367_),
	   .A (_net_7424) );
   NOR2_X1 g2636 (
	   .ZN (new_n9366_),
	   .A2 (n1993),
	   .A1 (new_n7739_) );
   NOR2_X1 g2635 (
	   .ZN (n3661),
	   .A2 (new_n7648_),
	   .A1 (new_n8543_) );
   CLKBUF_X1 g2634 (
	   .Z (n3658),
	   .A (net_6394) );
   CLKBUF_X1 g2633 (
	   .Z (n3655),
	   .A (net_6591) );
   CLKBUF_X1 g2632 (
	   .Z (n3651),
	   .A (net_7157) );
   OAI211_X1 g2631 (
	   .ZN (n3647),
	   .C2 (new_n7366_),
	   .C1 (new_n6852_),
	   .B (new_n9360_),
	   .A (new_n9359_) );
   NAND4_X1 g2630 (
	   .ZN (new_n9360_),
	   .A4 (_net_7718),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   NOR3_X1 g2629 (
	   .ZN (new_n9359_),
	   .A3 (new_n9358_),
	   .A2 (new_n9357_),
	   .A1 (new_n9356_1_) );
   AND3_X1 g2628 (
	   .ZN (new_n9358_),
	   .A3 (new_n7382_),
	   .A2 (net_257),
	   .A1 (new_n7380_) );
   NOR2_X1 g2627 (
	   .ZN (new_n9357_),
	   .A2 (new_n8505_),
	   .A1 (new_n7378_) );
   OAI22_X1 g2626 (
	   .ZN (new_n9356_1_),
	   .B2 (new_n9355_),
	   .B1 (new_n7938_),
	   .A2 (new_n9354_),
	   .A1 (new_n7936_) );
   INV_X1 g2625 (
	   .ZN (new_n9355_),
	   .A (net_183) );
   INV_X1 g2624 (
	   .ZN (new_n9354_),
	   .A (net_220) );
   NAND2_X1 g2623 (
	   .ZN (n3642),
	   .A2 (n4304),
	   .A1 (new_n7422_1_) );
   NOR2_X1 g2622 (
	   .ZN (n3638),
	   .A2 (new_n8193_),
	   .A1 (new_n9351_) );
   INV_X1 g2621 (
	   .ZN (new_n9351_),
	   .A (_net_190) );
   MUX2_X1 g2620 (
	   .Z (n3633),
	   .S (new_n7545_),
	   .B (_net_7665),
	   .A (new_n9349_) );
   OAI21_X1 g2619 (
	   .ZN (new_n9349_),
	   .B2 (new_n9348_1_),
	   .B1 (new_n7019_),
	   .A (new_n9347_) );
   INV_X1 g2618 (
	   .ZN (new_n9348_1_),
	   .A (net_371) );
   AOI22_X1 g2617 (
	   .ZN (new_n9347_),
	   .B2 (_net_292),
	   .B1 (net_383),
	   .A2 (_net_291),
	   .A1 (net_385) );
   OAI21_X1 g2616 (
	   .ZN (n3628),
	   .B2 (_net_7781),
	   .B1 (new_n9345_),
	   .A (new_n9343_1_) );
   NAND2_X1 g2615 (
	   .ZN (new_n9345_),
	   .A2 (new_n9342_),
	   .A1 (new_n9344_) );
   INV_X1 g2614 (
	   .ZN (new_n9344_),
	   .A (new_n9341_) );
   NAND3_X1 g2613 (
	   .ZN (new_n9343_1_),
	   .A3 (_net_7781),
	   .A2 (new_n9342_),
	   .A1 (new_n9341_) );
   INV_X1 g2612 (
	   .ZN (new_n9342_),
	   .A (_net_113) );
   NAND2_X1 g2611 (
	   .ZN (new_n9341_),
	   .A2 (new_n9340_),
	   .A1 (new_n7447_) );
   NAND3_X1 g2610 (
	   .ZN (new_n9340_),
	   .A3 (_net_7783),
	   .A2 (new_n9339_1_),
	   .A1 (new_n9338_) );
   INV_X1 g2609 (
	   .ZN (new_n9339_1_),
	   .A (_net_7782) );
   INV_X1 g2608 (
	   .ZN (new_n9338_),
	   .A (_net_7781) );
   CLKBUF_X1 g2607 (
	   .Z (n3623),
	   .A (_net_6124) );
   CLKBUF_X1 g2606 (
	   .Z (n3618),
	   .A (_net_7812) );
   MUX2_X1 g2605 (
	   .Z (n3614),
	   .S (new_n7437_1_),
	   .B (_net_5988),
	   .A (_net_7797) );
   NAND3_X1 g2604 (
	   .ZN (n3609),
	   .A3 (new_n9333_),
	   .A2 (new_n9332_),
	   .A1 (new_n9323_) );
   AOI22_X1 g2603 (
	   .ZN (new_n9333_),
	   .B2 (new_n7136_),
	   .B1 (net_6675),
	   .A2 (new_n7013_1_),
	   .A1 (new_n6975_) );
   AND3_X1 g2602 (
	   .ZN (new_n9332_),
	   .A3 (new_n9331_),
	   .A2 (new_n9330_1_),
	   .A1 (new_n9329_) );
   NAND2_X1 g2601 (
	   .ZN (new_n9331_),
	   .A2 (_net_6092),
	   .A1 (new_n6985_) );
   NAND2_X1 g2600 (
	   .ZN (new_n9330_1_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n8939_1_) );
   NAND2_X1 g2599 (
	   .ZN (new_n9329_),
	   .A2 (new_n6980_),
	   .A1 (new_n9328_) );
   NAND4_X1 g2598 (
	   .ZN (new_n9328_),
	   .A4 (new_n9327_),
	   .A3 (new_n9326_1_),
	   .A2 (new_n9325_),
	   .A1 (new_n9324_) );
   NAND3_X1 g2597 (
	   .ZN (new_n9327_),
	   .A3 (_net_6689),
	   .A2 (net_6663),
	   .A1 (_net_6688) );
   NAND3_X1 g2596 (
	   .ZN (new_n9326_1_),
	   .A3 (_net_6689),
	   .A2 (net_6631),
	   .A1 (new_n7004_) );
   NAND3_X1 g2595 (
	   .ZN (new_n9325_),
	   .A3 (_net_6688),
	   .A2 (net_6599),
	   .A1 (new_n7002_) );
   NAND2_X1 g2594 (
	   .ZN (new_n9324_),
	   .A2 (net_6567),
	   .A1 (new_n6973_) );
   AND3_X1 g2593 (
	   .ZN (new_n9323_),
	   .A3 (new_n9322_),
	   .A2 (new_n9321_1_),
	   .A1 (new_n9320_) );
   NAND4_X1 g2592 (
	   .ZN (new_n9322_),
	   .A4 (new_n6987_),
	   .A3 (net_6643),
	   .A2 (_net_6687),
	   .A1 (new_n7118_) );
   NAND4_X1 g2591 (
	   .ZN (new_n9321_1_),
	   .A4 (new_n6990_1_),
	   .A3 (_net_6687),
	   .A2 (net_6579),
	   .A1 (new_n7118_) );
   NAND4_X1 g2590 (
	   .ZN (new_n9320_),
	   .A4 (new_n6989_),
	   .A3 (net_6611),
	   .A2 (_net_6687),
	   .A1 (new_n7115_) );
   NOR2_X1 g2589 (
	   .ZN (n3604),
	   .A2 (new_n8000_),
	   .A1 (new_n7020_) );
   CLKBUF_X1 g2588 (
	   .Z (n3600),
	   .A (net_6583) );
   XNOR2_X1 g2587 (
	   .ZN (n3595),
	   .B (new_n9316_1_),
	   .A (new_n9315_) );
   NAND2_X1 g2586 (
	   .ZN (new_n9316_1_),
	   .A2 (net_6556),
	   .A1 (new_n6789_) );
   XNOR2_X1 g2585 (
	   .ZN (new_n9315_),
	   .B (_net_6557),
	   .A (_net_6554) );
   CLKBUF_X1 g2584 (
	   .Z (n3590),
	   .A (_net_7803) );
   CLKBUF_X1 g2583 (
	   .Z (n3587),
	   .A (net_6476) );
   NAND2_X1 g2582 (
	   .ZN (n3582),
	   .A2 (new_n9311_),
	   .A1 (new_n9310_) );
   AOI22_X1 g2581 (
	   .ZN (new_n9311_),
	   .B2 (_net_7577),
	   .B1 (new_n6755_),
	   .A2 (net_7609),
	   .A1 (new_n6743_) );
   AOI22_X1 g2580 (
	   .ZN (new_n9310_),
	   .B2 (net_7641),
	   .B1 (new_n8009_),
	   .A2 (new_n7970_1_),
	   .A1 (net_7673) );
   OAI21_X1 g2579 (
	   .ZN (n3577),
	   .B2 (new_n9308_),
	   .B1 (new_n9307_1_),
	   .A (new_n6963_) );
   NOR2_X1 g2578 (
	   .ZN (new_n9308_),
	   .A2 (_net_6408),
	   .A1 (new_n9305_) );
   NOR2_X1 g2577 (
	   .ZN (new_n9307_1_),
	   .A2 (new_n8185_),
	   .A1 (new_n9306_) );
   INV_X1 g2576 (
	   .ZN (new_n9306_),
	   .A (new_n9305_) );
   NOR2_X1 g2575 (
	   .ZN (new_n9305_),
	   .A2 (new_n9304_),
	   .A1 (new_n9303_) );
   INV_X1 g2574 (
	   .ZN (new_n9304_),
	   .A (_net_6407) );
   NAND3_X1 g2573 (
	   .ZN (new_n9303_),
	   .A3 (_net_6405),
	   .A2 (_net_6406),
	   .A1 (_net_6404) );
   MUX2_X1 g2572 (
	   .Z (n3572),
	   .S (new_n7285_),
	   .B (_net_7703),
	   .A (_net_7805) );
   AND2_X1 g2571 (
	   .ZN (n3567),
	   .A2 (net_378),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g2570 (
	   .Z (n3564),
	   .A (net_6873) );
   CLKBUF_X1 g2569 (
	   .Z (n3559),
	   .A (_net_7810) );
   CLKBUF_X1 g2568 (
	   .Z (n3555),
	   .A (net_6385) );
   AND2_X1 g2567 (
	   .ZN (n3551),
	   .A2 (_net_5983),
	   .A1 (_net_6039) );
   CLKBUF_X1 g2566 (
	   .Z (n3542),
	   .A (net_6885) );
   CLKBUF_X1 g2565 (
	   .Z (n3537),
	   .A (_net_6078) );
   CLKBUF_X1 g2564 (
	   .Z (n3532),
	   .A (net_6384) );
   CLKBUF_X1 g2563 (
	   .Z (n3528),
	   .A (_net_7815) );
   CLKBUF_X1 g2562 (
	   .Z (n3524),
	   .A (net_150) );
   CLKBUF_X1 g2561 (
	   .Z (n3520),
	   .A (_net_7800) );
   AOI21_X1 g2560 (
	   .ZN (n3516),
	   .B2 (new_n9288_),
	   .B1 (new_n6999_),
	   .A (new_n9289_) );
   OAI21_X1 g2559 (
	   .ZN (new_n9289_),
	   .B2 (new_n6999_),
	   .B1 (new_n9288_),
	   .A (_net_5995) );
   NAND2_X1 g2558 (
	   .ZN (new_n9288_),
	   .A2 (new_n6997_),
	   .A1 (new_n6982_1_) );
   CLKBUF_X1 g2557 (
	   .Z (n3511),
	   .A (_net_7793) );
   NAND3_X1 g2556 (
	   .ZN (n3507),
	   .A3 (new_n9285_),
	   .A2 (new_n9276_),
	   .A1 (new_n9270_) );
   AND3_X1 g2555 (
	   .ZN (new_n9285_),
	   .A3 (new_n9284_),
	   .A2 (new_n9283_),
	   .A1 (new_n9277_1_) );
   NAND2_X1 g2554 (
	   .ZN (new_n9284_),
	   .A2 (_net_6078),
	   .A1 (new_n6813_1_) );
   NAND2_X1 g2553 (
	   .ZN (new_n9283_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n9282_1_) );
   NAND4_X1 g2552 (
	   .ZN (new_n9282_1_),
	   .A4 (new_n9281_),
	   .A3 (new_n9280_),
	   .A2 (new_n9279_),
	   .A1 (new_n9278_) );
   NAND3_X1 g2551 (
	   .ZN (new_n9281_),
	   .A3 (net_6532),
	   .A2 (_net_6554),
	   .A1 (_net_6553) );
   NAND3_X1 g2550 (
	   .ZN (new_n9280_),
	   .A3 (_net_6554),
	   .A2 (net_6500),
	   .A1 (new_n6789_) );
   NAND3_X1 g2549 (
	   .ZN (new_n9279_),
	   .A3 (_net_6553),
	   .A2 (net_6468),
	   .A1 (new_n6787_) );
   NAND2_X1 g2548 (
	   .ZN (new_n9278_),
	   .A2 (net_6436),
	   .A1 (new_n6785_) );
   NAND2_X1 g2547 (
	   .ZN (new_n9277_1_),
	   .A2 (new_n7166_),
	   .A1 (new_n6792_) );
   AOI22_X1 g2546 (
	   .ZN (new_n9276_),
	   .B2 (new_n9275_),
	   .B1 (new_n6784_),
	   .A2 (new_n6779_1_),
	   .A1 (net_6546) );
   NAND4_X1 g2545 (
	   .ZN (new_n9275_),
	   .A4 (new_n9274_),
	   .A3 (new_n9273_),
	   .A2 (new_n9272_1_),
	   .A1 (new_n9271_) );
   NAND3_X1 g2544 (
	   .ZN (new_n9274_),
	   .A3 (_net_6554),
	   .A2 (net_6530),
	   .A1 (_net_6553) );
   NAND3_X1 g2543 (
	   .ZN (new_n9273_),
	   .A3 (_net_6554),
	   .A2 (net_6498),
	   .A1 (new_n6789_) );
   NAND3_X1 g2542 (
	   .ZN (new_n9272_1_),
	   .A3 (net_6466),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   NAND2_X1 g2541 (
	   .ZN (new_n9271_),
	   .A2 (net_6434),
	   .A1 (new_n6785_) );
   AND3_X1 g2540 (
	   .ZN (new_n9270_),
	   .A3 (new_n9269_),
	   .A2 (new_n9268_),
	   .A1 (new_n9267_1_) );
   NAND4_X1 g2539 (
	   .ZN (new_n9269_),
	   .A4 (new_n6775_),
	   .A3 (_net_6552),
	   .A2 (net_6514),
	   .A1 (new_n6772_) );
   NAND4_X1 g2538 (
	   .ZN (new_n9268_),
	   .A4 (new_n6770_1_),
	   .A3 (_net_6552),
	   .A2 (net_6450),
	   .A1 (new_n6772_) );
   NAND4_X1 g2537 (
	   .ZN (new_n9267_1_),
	   .A4 (new_n6767_),
	   .A3 (_net_6552),
	   .A2 (net_6482),
	   .A1 (new_n6764_) );
   CLKBUF_X1 g2536 (
	   .Z (n3502),
	   .A (_net_263) );
   CLKBUF_X1 g2535 (
	   .Z (n3497),
	   .A (_net_7803) );
   CLKBUF_X1 g2534 (
	   .Z (n3494),
	   .A (net_7241) );
   OAI21_X1 g2533 (
	   .ZN (n3489),
	   .B2 (new_n7111_1_),
	   .B1 (new_n9262_),
	   .A (new_n9261_) );
   INV_X1 g2532 (
	   .ZN (new_n9262_),
	   .A (_net_7362) );
   NAND2_X1 g2531 (
	   .ZN (new_n9261_),
	   .A2 (new_n7321_1_),
	   .A1 (new_n7101_) );
   AND2_X1 g2530 (
	   .ZN (n3484),
	   .A2 (_net_6289),
	   .A1 (new_n7239_) );
   CLKBUF_X1 g2529 (
	   .Z (n3479),
	   .A (_net_6136) );
   NAND4_X1 g2528 (
	   .ZN (n3474),
	   .A4 (new_n9257_),
	   .A3 (new_n9256_),
	   .A2 (new_n9254_1_),
	   .A1 (new_n9250_1_) );
   AOI22_X1 g2527 (
	   .ZN (new_n9257_),
	   .B2 (_net_6130),
	   .B1 (new_n6869_),
	   .A2 (new_n6854_),
	   .A1 (new_n8502_) );
   NAND2_X1 g2526 (
	   .ZN (new_n9256_),
	   .A2 (new_n9184_),
	   .A1 (new_n9255_) );
   NOR2_X1 g2525 (
	   .ZN (new_n9255_),
	   .A2 (new_n8591_),
	   .A1 (new_n6877_) );
   NAND2_X1 g2524 (
	   .ZN (new_n9254_1_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n9253_) );
   NAND2_X1 g2523 (
	   .ZN (new_n9253_),
	   .A2 (new_n9252_),
	   .A1 (new_n9251_) );
   AOI22_X1 g2522 (
	   .ZN (new_n9252_),
	   .B2 (net_6833),
	   .B1 (new_n6844_),
	   .A2 (net_6865),
	   .A1 (new_n6832_) );
   AOI22_X1 g2521 (
	   .ZN (new_n9251_),
	   .B2 (net_6929),
	   .B1 (new_n6873_),
	   .A2 (new_n6840_1_),
	   .A1 (net_6897) );
   NAND2_X1 g2520 (
	   .ZN (new_n9250_1_),
	   .A2 (new_n6879_),
	   .A1 (new_n9249_) );
   NAND2_X1 g2519 (
	   .ZN (new_n9249_),
	   .A2 (new_n9248_),
	   .A1 (new_n9247_) );
   AOI22_X1 g2518 (
	   .ZN (new_n9248_),
	   .B2 (net_6831),
	   .B1 (new_n6836_1_),
	   .A2 (net_6863),
	   .A1 (new_n6833_) );
   AOI22_X1 g2517 (
	   .ZN (new_n9247_),
	   .B2 (net_6927),
	   .B1 (new_n6873_),
	   .A2 (new_n6841_),
	   .A1 (net_6895) );
   CLKBUF_X1 g2516 (
	   .Z (n3469),
	   .A (_net_7811) );
   XNOR2_X1 g2515 (
	   .ZN (n3464),
	   .B (_net_7382),
	   .A (net_7378) );
   NAND3_X1 g2514 (
	   .ZN (n3459),
	   .A3 (new_n9243_),
	   .A2 (new_n9239_),
	   .A1 (new_n9233_1_) );
   AND3_X1 g2513 (
	   .ZN (new_n9243_),
	   .A3 (new_n9242_1_),
	   .A2 (new_n9241_),
	   .A1 (new_n9240_) );
   NAND2_X1 g2512 (
	   .ZN (new_n9242_1_),
	   .A2 (_net_6075),
	   .A1 (new_n6813_1_) );
   NAND2_X1 g2511 (
	   .ZN (new_n9241_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n8079_) );
   NAND2_X1 g2510 (
	   .ZN (new_n9240_),
	   .A2 (new_n7166_),
	   .A1 (new_n7159_) );
   AOI22_X1 g2509 (
	   .ZN (new_n9239_),
	   .B2 (new_n9238_1_),
	   .B1 (new_n6784_),
	   .A2 (new_n6779_1_),
	   .A1 (net_6543) );
   NAND4_X1 g2508 (
	   .ZN (new_n9238_1_),
	   .A4 (new_n9237_),
	   .A3 (new_n9236_),
	   .A2 (new_n9235_),
	   .A1 (new_n9234_) );
   NAND3_X1 g2507 (
	   .ZN (new_n9237_),
	   .A3 (net_6527),
	   .A2 (_net_6554),
	   .A1 (_net_6553) );
   NAND3_X1 g2506 (
	   .ZN (new_n9236_),
	   .A3 (_net_6554),
	   .A2 (net_6495),
	   .A1 (new_n6789_) );
   NAND3_X1 g2505 (
	   .ZN (new_n9235_),
	   .A3 (net_6463),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   NAND2_X1 g2504 (
	   .ZN (new_n9234_),
	   .A2 (net_6431),
	   .A1 (new_n6785_) );
   AND3_X1 g2503 (
	   .ZN (new_n9233_1_),
	   .A3 (new_n9232_),
	   .A2 (new_n9231_),
	   .A1 (new_n9230_) );
   NAND4_X1 g2502 (
	   .ZN (new_n9232_),
	   .A4 (new_n6775_),
	   .A3 (_net_6552),
	   .A2 (net_6511),
	   .A1 (new_n6772_) );
   NAND4_X1 g2501 (
	   .ZN (new_n9231_),
	   .A4 (new_n6770_1_),
	   .A3 (_net_6552),
	   .A2 (net_6447),
	   .A1 (new_n6772_) );
   NAND4_X1 g2500 (
	   .ZN (new_n9230_),
	   .A4 (new_n6767_),
	   .A3 (_net_6552),
	   .A2 (net_6479),
	   .A1 (new_n6764_) );
   NAND3_X1 g2499 (
	   .ZN (n3455),
	   .A3 (new_n9228_1_),
	   .A2 (new_n9227_),
	   .A1 (new_n9219_) );
   OR2_X1 g2498 (
	   .ZN (new_n9228_1_),
	   .A2 (new_n6811_),
	   .A1 (new_n7365_) );
   NOR3_X1 g2497 (
	   .ZN (new_n9227_),
	   .A3 (new_n9226_),
	   .A2 (new_n9222_),
	   .A1 (new_n9220_1_) );
   NAND3_X1 g2496 (
	   .ZN (new_n9226_),
	   .A3 (new_n9225_1_),
	   .A2 (new_n9224_),
	   .A1 (new_n9223_) );
   NAND4_X1 g2495 (
	   .ZN (new_n9225_1_),
	   .A4 (net_156),
	   .A3 (x1231),
	   .A2 (new_n7394_),
	   .A1 (new_n7393_) );
   NAND3_X1 g2494 (
	   .ZN (new_n9224_),
	   .A3 (_net_193),
	   .A2 (new_n7388_),
	   .A1 (new_n7387_) );
   NAND3_X1 g2493 (
	   .ZN (new_n9223_),
	   .A3 (net_230),
	   .A2 (new_n7383_),
	   .A1 (new_n7380_) );
   OAI22_X1 g2492 (
	   .ZN (new_n9222_),
	   .B2 (new_n7378_),
	   .B1 (new_n8540_1_),
	   .A2 (new_n9221_),
	   .A1 (new_n7374_) );
   INV_X1 g2491 (
	   .ZN (new_n9221_),
	   .A (_net_114) );
   AND4_X1 g2490 (
	   .ZN (new_n9220_1_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7369_),
	   .A1 (_net_6028) );
   NOR2_X1 g2489 (
	   .ZN (new_n9219_),
	   .A2 (new_n9218_),
	   .A1 (new_n9217_) );
   NOR2_X1 g2488 (
	   .ZN (new_n9218_),
	   .A2 (new_n8193_),
	   .A1 (new_n7362_) );
   NOR2_X1 g2487 (
	   .ZN (new_n9217_),
	   .A2 (new_n9216_),
	   .A1 (new_n9215_1_) );
   INV_X1 g2486 (
	   .ZN (new_n9216_),
	   .A (net_7691) );
   NAND4_X1 g2485 (
	   .ZN (new_n9215_1_),
	   .A4 (new_n7360_),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7357_) );
   CLKBUF_X1 g2484 (
	   .Z (n3450),
	   .A (_net_6173) );
   CLKBUF_X1 g2483 (
	   .Z (n3445),
	   .A (net_6389) );
   OAI221_X1 g2482 (
	   .ZN (n3440),
	   .C2 (new_n7306_),
	   .C1 (new_n9211_1_),
	   .B2 (new_n7303_),
	   .B1 (new_n8282_),
	   .A (new_n9210_) );
   INV_X1 g2481 (
	   .ZN (new_n9211_1_),
	   .A (_net_7515) );
   AOI22_X1 g2480 (
	   .ZN (new_n9210_),
	   .B2 (_net_7419),
	   .B1 (new_n9203_),
	   .A2 (_net_7451),
	   .A1 (new_n8694_1_) );
   CLKBUF_X1 g2479 (
	   .Z (n3436),
	   .A (net_7120) );
   NAND2_X1 g2478 (
	   .ZN (n3431),
	   .A2 (n4304),
	   .A1 (new_n7422_1_) );
   MUX2_X1 g2477 (
	   .Z (n3427),
	   .S (new_n7504_),
	   .B (_net_7618),
	   .A (new_n8114_) );
   OAI221_X1 g2476 (
	   .ZN (n3422),
	   .C2 (new_n7303_),
	   .C1 (new_n9205_),
	   .B2 (new_n7306_),
	   .B1 (new_n8861_),
	   .A (new_n9204_) );
   INV_X1 g2475 (
	   .ZN (new_n9205_),
	   .A (_net_7469) );
   AOI22_X1 g2474 (
	   .ZN (new_n9204_),
	   .B2 (_net_7405),
	   .B1 (new_n9203_),
	   .A2 (_net_7437),
	   .A1 (new_n8694_1_) );
   BUF_X4 g2473 (
	   .Z (new_n9203_),
	   .A (new_n7297_1_) );
   CLKBUF_X1 g2472 (
	   .Z (n3418),
	   .A (net_7248) );
   CLKBUF_X1 g2471 (
	   .Z (n3413),
	   .A (net_148) );
   CLKBUF_X1 g2470 (
	   .Z (n3408),
	   .A (_net_7820) );
   CLKBUF_X1 g2469 (
	   .Z (n3404),
	   .A (net_6386) );
   MUX2_X1 g2468 (
	   .Z (n3400),
	   .S (new_n7504_),
	   .B (_net_7619),
	   .A (new_n9197_) );
   OAI21_X1 g2467 (
	   .ZN (new_n9197_),
	   .B2 (new_n9196_1_),
	   .B1 (new_n7019_),
	   .A (new_n9195_) );
   INV_X1 g2466 (
	   .ZN (new_n9196_1_),
	   .A (net_7539) );
   AOI22_X1 g2465 (
	   .ZN (new_n9195_),
	   .B2 (_net_292),
	   .B1 (net_369),
	   .A2 (_net_291),
	   .A1 (net_371) );
   NAND3_X1 g2464 (
	   .ZN (n3395),
	   .A3 (new_n9193_),
	   .A2 (new_n9187_1_),
	   .A1 (new_n9173_1_) );
   AOI22_X1 g2463 (
	   .ZN (new_n9193_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6955),
	   .A2 (new_n9192_1_),
	   .A1 (new_n6879_) );
   NAND4_X1 g2462 (
	   .ZN (new_n9192_1_),
	   .A4 (new_n9191_),
	   .A3 (new_n9190_),
	   .A2 (new_n9189_),
	   .A1 (new_n9188_) );
   NAND3_X1 g2461 (
	   .ZN (new_n9191_),
	   .A3 (_net_6958),
	   .A2 (_net_6959),
	   .A1 (net_6939) );
   NAND3_X1 g2460 (
	   .ZN (new_n9190_),
	   .A3 (_net_6959),
	   .A2 (net_6907),
	   .A1 (new_n6848_) );
   NAND3_X1 g2459 (
	   .ZN (new_n9189_),
	   .A3 (_net_6958),
	   .A2 (net_6875),
	   .A1 (new_n6846_) );
   NAND2_X1 g2458 (
	   .ZN (new_n9188_),
	   .A2 (net_6843),
	   .A1 (new_n6844_) );
   AND3_X1 g2457 (
	   .ZN (new_n9187_1_),
	   .A3 (new_n9186_),
	   .A2 (new_n9185_),
	   .A1 (new_n9179_) );
   NAND2_X1 g2456 (
	   .ZN (new_n9186_),
	   .A2 (_net_6142),
	   .A1 (new_n6869_) );
   NAND2_X1 g2455 (
	   .ZN (new_n9185_),
	   .A2 (new_n6853_),
	   .A1 (new_n9184_) );
   NAND4_X1 g2454 (
	   .ZN (new_n9184_),
	   .A4 (new_n9183_),
	   .A3 (new_n9182_1_),
	   .A2 (new_n9181_),
	   .A1 (new_n9180_) );
   NAND3_X1 g2453 (
	   .ZN (new_n9183_),
	   .A3 (net_6943),
	   .A2 (_net_6958),
	   .A1 (_net_6959) );
   NAND3_X1 g2452 (
	   .ZN (new_n9182_1_),
	   .A3 (net_6911),
	   .A2 (_net_6959),
	   .A1 (new_n6848_) );
   NAND3_X1 g2451 (
	   .ZN (new_n9181_),
	   .A3 (net_6879),
	   .A2 (_net_6958),
	   .A1 (new_n6846_) );
   NAND2_X1 g2450 (
	   .ZN (new_n9180_),
	   .A2 (net_6847),
	   .A1 (new_n6844_) );
   NAND2_X1 g2449 (
	   .ZN (new_n9179_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n9178_1_) );
   NAND4_X1 g2448 (
	   .ZN (new_n9178_1_),
	   .A4 (new_n9177_),
	   .A3 (new_n9176_),
	   .A2 (new_n9175_),
	   .A1 (new_n9174_) );
   NAND3_X1 g2447 (
	   .ZN (new_n9177_),
	   .A3 (_net_6958),
	   .A2 (_net_6959),
	   .A1 (net_6941) );
   NAND3_X1 g2446 (
	   .ZN (new_n9176_),
	   .A3 (_net_6959),
	   .A2 (net_6909),
	   .A1 (new_n6848_) );
   NAND3_X1 g2445 (
	   .ZN (new_n9175_),
	   .A3 (_net_6958),
	   .A2 (net_6877),
	   .A1 (new_n6846_) );
   NAND2_X1 g2444 (
	   .ZN (new_n9174_),
	   .A2 (net_6845),
	   .A1 (new_n6844_) );
   AND3_X1 g2443 (
	   .ZN (new_n9173_1_),
	   .A3 (new_n9172_),
	   .A2 (new_n9171_),
	   .A1 (new_n9170_) );
   NAND4_X1 g2442 (
	   .ZN (new_n9172_),
	   .A4 (new_n6841_),
	   .A3 (_net_6957),
	   .A2 (net_6923),
	   .A1 (new_n6838_) );
   NAND4_X1 g2441 (
	   .ZN (new_n9171_),
	   .A4 (new_n6836_1_),
	   .A3 (_net_6957),
	   .A2 (net_6859),
	   .A1 (new_n6838_) );
   NAND4_X1 g2440 (
	   .ZN (new_n9170_),
	   .A4 (new_n6833_),
	   .A3 (net_6891),
	   .A2 (_net_6957),
	   .A1 (new_n6830_) );
   CLKBUF_X1 g2439 (
	   .Z (n3390),
	   .A (x1424) );
   CLKBUF_X1 g2438 (
	   .Z (n3386),
	   .A (net_7807) );
   CLKBUF_X1 g2437 (
	   .Z (n3383),
	   .A (net_6485) );
   CLKBUF_X1 g2436 (
	   .Z (n3379),
	   .A (net_6698) );
   NOR2_X1 g2435 (
	   .ZN (n3374),
	   .A2 (new_n7275_1_),
	   .A1 (new_n8543_) );
   NOR4_X1 g2434 (
	   .ZN (n3370),
	   .A4 (new_n9163_),
	   .A3 (new_n9162_),
	   .A2 (new_n9161_),
	   .A1 (new_n9158_) );
   NOR2_X1 g2433 (
	   .ZN (new_n9163_),
	   .A2 (_net_7232),
	   .A1 (new_n8383_) );
   NOR2_X1 g2432 (
	   .ZN (new_n9162_),
	   .A2 (new_n7843_),
	   .A1 (new_n9155_) );
   NAND2_X1 g2431 (
	   .ZN (new_n9161_),
	   .A2 (new_n9160_1_),
	   .A1 (new_n9159_) );
   NAND2_X1 g2430 (
	   .ZN (new_n9160_1_),
	   .A2 (_net_7232),
	   .A1 (new_n8383_) );
   OAI21_X1 g2429 (
	   .ZN (new_n9159_),
	   .B2 (new_n7810_1_),
	   .B1 (n4276),
	   .A (_net_7227) );
   OAI21_X1 g2428 (
	   .ZN (new_n9158_),
	   .B2 (n4276),
	   .B1 (_net_7227),
	   .A (new_n9156_1_) );
   XNOR2_X1 g2427 (
	   .ZN (n4276),
	   .B (_net_7228),
	   .A (net_7231) );
   NAND2_X1 g2426 (
	   .ZN (new_n9156_1_),
	   .A2 (new_n7843_),
	   .A1 (new_n9155_) );
   XOR2_X1 g2425 (
	   .Z (new_n9155_),
	   .B (_net_7230),
	   .A (_net_7233) );
   CLKBUF_X1 g2424 (
	   .Z (n3365),
	   .A (_net_7821) );
   CLKBUF_X1 g2423 (
	   .Z (n3361),
	   .A (_net_6071) );
   MUX2_X1 g2422 (
	   .Z (n3356),
	   .S (new_n7609_),
	   .B (_net_7583),
	   .A (n5628) );
   NOR2_X1 g2421 (
	   .ZN (n5628),
	   .A2 (new_n7214_),
	   .A1 (new_n7020_) );
   NAND3_X1 g2420 (
	   .ZN (n3352),
	   .A3 (new_n9149_),
	   .A2 (new_n9148_),
	   .A1 (new_n9139_) );
   NAND4_X1 g2419 (
	   .ZN (new_n9149_),
	   .A4 (_net_7700),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR3_X1 g2418 (
	   .ZN (new_n9148_),
	   .A3 (new_n9147_),
	   .A2 (new_n9143_1_),
	   .A1 (new_n9140_) );
   NAND3_X1 g2417 (
	   .ZN (new_n9147_),
	   .A3 (new_n9146_1_),
	   .A2 (new_n9145_),
	   .A1 (new_n9144_) );
   NAND4_X1 g2416 (
	   .ZN (new_n9146_1_),
	   .A4 (net_165),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g2415 (
	   .ZN (new_n9145_),
	   .A3 (net_202),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g2414 (
	   .ZN (new_n9144_),
	   .A3 (net_239),
	   .A2 (new_n7383_),
	   .A1 (new_n7380_) );
   OAI22_X1 g2413 (
	   .ZN (new_n9143_1_),
	   .B2 (new_n7378_),
	   .B1 (new_n9142_),
	   .A2 (new_n9141_),
	   .A1 (new_n7374_) );
   INV_X1 g2412 (
	   .ZN (new_n9142_),
	   .A (_net_7729) );
   INV_X1 g2411 (
	   .ZN (new_n9141_),
	   .A (_net_123) );
   AND4_X1 g2410 (
	   .ZN (new_n9140_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7369_),
	   .A1 (_net_6040) );
   NOR2_X1 g2409 (
	   .ZN (new_n9139_),
	   .A2 (new_n9138_1_),
	   .A1 (new_n9136_) );
   NOR2_X1 g2408 (
	   .ZN (new_n9138_1_),
	   .A2 (new_n9137_),
	   .A1 (new_n7366_) );
   INV_X1 g2407 (
	   .ZN (new_n9137_),
	   .A (_net_5996) );
   NOR2_X1 g2406 (
	   .ZN (new_n9136_),
	   .A2 (new_n9135_),
	   .A1 (new_n7362_) );
   INV_X1 g2405 (
	   .ZN (new_n9135_),
	   .A (_net_279) );
   CLKBUF_X1 g2404 (
	   .Z (n3348),
	   .A (net_7140) );
   CLKBUF_X1 g2403 (
	   .Z (n3343),
	   .A (_net_6063) );
   MUX2_X1 g2402 (
	   .Z (n3338),
	   .S (new_n6823_),
	   .B (_net_6041),
	   .A (_net_7803) );
   NOR2_X1 g2401 (
	   .ZN (n3333),
	   .A2 (new_n7334_),
	   .A1 (new_n8675_) );
   CLKBUF_X1 g2400 (
	   .Z (n3330),
	   .A (net_6868) );
   AND2_X1 g2399 (
	   .ZN (n3325),
	   .A2 (net_342),
	   .A1 (new_n7102_1_) );
   NAND4_X1 g2398 (
	   .ZN (n3322),
	   .A4 (new_n9127_),
	   .A3 (new_n9126_),
	   .A2 (new_n9125_),
	   .A1 (new_n9124_1_) );
   NAND4_X1 g2397 (
	   .ZN (new_n9127_),
	   .A4 (new_n7364_),
	   .A3 (_net_6002),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   NAND4_X1 g2396 (
	   .ZN (new_n9126_),
	   .A4 (_net_7706),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   NAND4_X1 g2395 (
	   .ZN (new_n9125_),
	   .A4 (net_285),
	   .A3 (x1286),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR2_X1 g2394 (
	   .ZN (new_n9124_1_),
	   .A2 (new_n9123_),
	   .A1 (new_n9118_) );
   NAND4_X1 g2393 (
	   .ZN (new_n9123_),
	   .A4 (new_n9122_),
	   .A3 (new_n9121_),
	   .A2 (new_n9120_1_),
	   .A1 (new_n9119_) );
   NAND4_X1 g2392 (
	   .ZN (new_n9122_),
	   .A4 (net_171),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g2391 (
	   .ZN (new_n9121_),
	   .A3 (net_208),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g2390 (
	   .ZN (new_n9120_1_),
	   .A3 (net_245),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   NAND4_X1 g2389 (
	   .ZN (new_n9119_),
	   .A4 (_net_7735),
	   .A3 (x1286),
	   .A2 (x1261),
	   .A1 (new_n7370_) );
   NAND2_X1 g2388 (
	   .ZN (new_n9118_),
	   .A2 (new_n9117_),
	   .A1 (new_n9116_) );
   NAND4_X1 g2387 (
	   .ZN (new_n9117_),
	   .A4 (new_n7354_1_),
	   .A3 (_net_129),
	   .A2 (x1261),
	   .A1 (new_n7370_) );
   NAND4_X1 g2386 (
	   .ZN (new_n9116_),
	   .A4 (new_n7371_),
	   .A3 (new_n7370_),
	   .A2 (net_6046),
	   .A1 (new_n7369_) );
   CLKBUF_X1 g2385 (
	   .Z (n3318),
	   .A (net_6883) );
   NAND4_X1 g2384 (
	   .ZN (n3313),
	   .A4 (new_n9113_),
	   .A3 (new_n9112_),
	   .A2 (new_n9111_),
	   .A1 (new_n9110_1_) );
   AOI22_X1 g2383 (
	   .ZN (new_n9113_),
	   .B2 (_net_6171),
	   .B1 (new_n7694_),
	   .A2 (new_n7690_),
	   .A1 (new_n9057_1_) );
   NAND2_X1 g2382 (
	   .ZN (new_n9112_),
	   .A2 (new_n7701_),
	   .A1 (new_n8547_) );
   NAND2_X1 g2381 (
	   .ZN (new_n9111_),
	   .A2 (new_n7837_),
	   .A1 (new_n7685_) );
   NAND2_X1 g2380 (
	   .ZN (new_n9110_1_),
	   .A2 (new_n9109_),
	   .A1 (new_n8026_) );
   NAND4_X1 g2379 (
	   .ZN (new_n9109_),
	   .A4 (new_n9108_),
	   .A3 (new_n9107_),
	   .A2 (new_n9106_1_),
	   .A1 (new_n9105_) );
   NAND3_X1 g2378 (
	   .ZN (new_n9108_),
	   .A3 (net_7214),
	   .A2 (_net_7228),
	   .A1 (_net_7229) );
   NAND3_X1 g2377 (
	   .ZN (new_n9107_),
	   .A3 (_net_7229),
	   .A2 (net_7182),
	   .A1 (new_n7823_) );
   NAND3_X1 g2376 (
	   .ZN (new_n9106_1_),
	   .A3 (_net_7228),
	   .A2 (net_7150),
	   .A1 (new_n7821_) );
   NAND2_X1 g2375 (
	   .ZN (new_n9105_),
	   .A2 (net_7118),
	   .A1 (new_n7819_) );
   OAI21_X1 g2374 (
	   .ZN (n3308),
	   .B2 (new_n6957_1_),
	   .B1 (new_n9103_),
	   .A (new_n9102_) );
   INV_X1 g2373 (
	   .ZN (new_n9103_),
	   .A (_net_7266) );
   NAND2_X1 g2372 (
	   .ZN (new_n9102_),
	   .A2 (new_n7321_1_),
	   .A1 (new_n6949_) );
   CLKBUF_X1 g2371 (
	   .Z (n3303),
	   .A (_net_7809) );
   CLKBUF_X1 g2370 (
	   .Z (n3299),
	   .A (_net_7793) );
   NAND3_X1 g2369 (
	   .ZN (n3294),
	   .A3 (new_n9098_),
	   .A2 (new_n9084_),
	   .A1 (new_n9083_) );
   AND3_X1 g2368 (
	   .ZN (new_n9098_),
	   .A3 (new_n9097_),
	   .A2 (new_n9096_1_),
	   .A1 (new_n9090_) );
   NAND2_X1 g2367 (
	   .ZN (new_n9097_),
	   .A2 (_net_6083),
	   .A1 (new_n6813_1_) );
   NAND2_X1 g2366 (
	   .ZN (new_n9096_1_),
	   .A2 (new_n6809_1_),
	   .A1 (new_n9095_) );
   NAND4_X1 g2365 (
	   .ZN (new_n9095_),
	   .A4 (new_n9094_),
	   .A3 (new_n9093_),
	   .A2 (new_n9092_),
	   .A1 (new_n9091_1_) );
   NAND3_X1 g2364 (
	   .ZN (new_n9094_),
	   .A3 (_net_6554),
	   .A2 (_net_6553),
	   .A1 (net_6539) );
   NAND3_X1 g2363 (
	   .ZN (new_n9093_),
	   .A3 (net_6507),
	   .A2 (_net_6554),
	   .A1 (new_n6789_) );
   NAND3_X1 g2362 (
	   .ZN (new_n9092_),
	   .A3 (net_6475),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   NAND2_X1 g2361 (
	   .ZN (new_n9091_1_),
	   .A2 (net_6443),
	   .A1 (new_n6785_) );
   NAND2_X1 g2360 (
	   .ZN (new_n9090_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n9089_) );
   NAND4_X1 g2359 (
	   .ZN (new_n9089_),
	   .A4 (new_n9088_),
	   .A3 (new_n9087_),
	   .A2 (new_n9086_1_),
	   .A1 (new_n9085_) );
   NAND3_X1 g2358 (
	   .ZN (new_n9088_),
	   .A3 (_net_6554),
	   .A2 (_net_6553),
	   .A1 (net_6537) );
   NAND3_X1 g2357 (
	   .ZN (new_n9087_),
	   .A3 (_net_6554),
	   .A2 (net_6505),
	   .A1 (new_n6789_) );
   NAND3_X1 g2356 (
	   .ZN (new_n9086_1_),
	   .A3 (net_6473),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   NAND2_X1 g2355 (
	   .ZN (new_n9085_),
	   .A2 (net_6441),
	   .A1 (new_n6785_) );
   AOI22_X1 g2354 (
	   .ZN (new_n9084_),
	   .B2 (new_n7165_),
	   .B1 (new_n6784_),
	   .A2 (new_n6779_1_),
	   .A1 (net_6551) );
   AND3_X1 g2353 (
	   .ZN (new_n9083_),
	   .A3 (new_n9082_1_),
	   .A2 (new_n9081_),
	   .A1 (new_n9080_) );
   NAND4_X1 g2352 (
	   .ZN (new_n9082_1_),
	   .A4 (new_n6775_),
	   .A3 (_net_6552),
	   .A2 (net_6519),
	   .A1 (new_n6772_) );
   NAND4_X1 g2351 (
	   .ZN (new_n9081_),
	   .A4 (new_n6770_1_),
	   .A3 (net_6455),
	   .A2 (_net_6552),
	   .A1 (new_n6772_) );
   NAND4_X1 g2350 (
	   .ZN (new_n9080_),
	   .A4 (new_n6767_),
	   .A3 (_net_6552),
	   .A2 (net_6487),
	   .A1 (new_n6764_) );
   CLKBUF_X1 g2349 (
	   .Z (n3290),
	   .A (net_7710) );
   AND2_X1 g2348 (
	   .ZN (n3285),
	   .A2 (_net_6203),
	   .A1 (new_n7239_) );
   CLKBUF_X1 g2347 (
	   .Z (n3280),
	   .A (_net_7795) );
   NOR2_X1 g2346 (
	   .ZN (n3276),
	   .A2 (new_n6933_),
	   .A1 (new_n8543_) );
   CLKBUF_X1 g2345 (
	   .Z (n3272),
	   .A (net_7799) );
   NAND3_X1 g2344 (
	   .ZN (n3268),
	   .A3 (new_n9073_),
	   .A2 (new_n9072_),
	   .A1 (new_n9068_) );
   AOI22_X1 g2343 (
	   .ZN (new_n9073_),
	   .B2 (new_n7136_),
	   .B1 (net_6685),
	   .A2 (new_n7126_),
	   .A1 (new_n7013_1_) );
   AND3_X1 g2342 (
	   .ZN (new_n9072_),
	   .A3 (new_n9071_),
	   .A2 (new_n9070_),
	   .A1 (new_n9069_1_) );
   NAND2_X1 g2341 (
	   .ZN (new_n9071_),
	   .A2 (_net_6102),
	   .A1 (new_n6985_) );
   NAND2_X1 g2340 (
	   .ZN (new_n9070_),
	   .A2 (new_n6979_),
	   .A1 (new_n8933_) );
   NAND2_X1 g2339 (
	   .ZN (new_n9069_1_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n7007_) );
   AND3_X1 g2338 (
	   .ZN (new_n9068_),
	   .A3 (new_n9067_),
	   .A2 (new_n9066_),
	   .A1 (new_n9065_1_) );
   NAND4_X1 g2337 (
	   .ZN (new_n9067_),
	   .A4 (new_n6987_),
	   .A3 (_net_6687),
	   .A2 (net_6653),
	   .A1 (new_n7118_) );
   NAND4_X1 g2336 (
	   .ZN (new_n9066_),
	   .A4 (new_n6990_1_),
	   .A3 (net_6589),
	   .A2 (_net_6687),
	   .A1 (new_n7118_) );
   NAND4_X1 g2335 (
	   .ZN (new_n9065_1_),
	   .A4 (new_n6989_),
	   .A3 (net_6621),
	   .A2 (_net_6687),
	   .A1 (new_n7115_) );
   MUX2_X1 g2334 (
	   .Z (n3263),
	   .S (_net_154),
	   .B (net_312),
	   .A (_net_116) );
   CLKBUF_X1 g2333 (
	   .Z (n3258),
	   .A (x1366) );
   MUX2_X1 g2332 (
	   .Z (n3254),
	   .S (new_n7538_),
	   .B (_net_272),
	   .A (_net_7798) );
   CLKBUF_X1 g2331 (
	   .Z (n3249),
	   .A (_net_6083) );
   CLKBUF_X1 g2330 (
	   .Z (n3244),
	   .A (_net_7822) );
   NAND3_X1 g2329 (
	   .ZN (n3240),
	   .A3 (new_n9058_),
	   .A2 (new_n9052_1_),
	   .A1 (new_n9048_) );
   AOI22_X1 g2328 (
	   .ZN (new_n9058_),
	   .B2 (net_7218),
	   .B1 (new_n7844_),
	   .A2 (new_n9057_1_),
	   .A1 (new_n7837_) );
   NAND4_X1 g2327 (
	   .ZN (new_n9057_1_),
	   .A4 (new_n9056_),
	   .A3 (new_n9055_),
	   .A2 (new_n9054_),
	   .A1 (new_n9053_) );
   NAND3_X1 g2326 (
	   .ZN (new_n9056_),
	   .A3 (_net_7228),
	   .A2 (net_7202),
	   .A1 (_net_7229) );
   NAND3_X1 g2325 (
	   .ZN (new_n9055_),
	   .A3 (_net_7229),
	   .A2 (net_7170),
	   .A1 (new_n7823_) );
   NAND3_X1 g2324 (
	   .ZN (new_n9054_),
	   .A3 (net_7138),
	   .A2 (_net_7228),
	   .A1 (new_n7821_) );
   NAND2_X1 g2323 (
	   .ZN (new_n9053_),
	   .A2 (net_7106),
	   .A1 (new_n7819_) );
   AND3_X1 g2322 (
	   .ZN (new_n9052_1_),
	   .A3 (new_n9051_),
	   .A2 (new_n9050_),
	   .A1 (new_n9049_) );
   NAND2_X1 g2321 (
	   .ZN (new_n9051_),
	   .A2 (_net_6175),
	   .A1 (new_n7694_) );
   NAND2_X1 g2320 (
	   .ZN (new_n9050_),
	   .A2 (new_n7701_),
	   .A1 (new_n8376_) );
   NAND2_X1 g2319 (
	   .ZN (new_n9049_),
	   .A2 (new_n7690_),
	   .A1 (new_n8368_) );
   AND3_X1 g2318 (
	   .ZN (new_n9048_),
	   .A3 (new_n9047_1_),
	   .A2 (new_n9046_),
	   .A1 (new_n9045_) );
   NAND4_X1 g2317 (
	   .ZN (new_n9047_1_),
	   .A4 (new_n7678_),
	   .A3 (net_7186),
	   .A2 (_net_7227),
	   .A1 (new_n7816_) );
   NAND4_X1 g2316 (
	   .ZN (new_n9046_),
	   .A4 (new_n7683_),
	   .A3 (net_7122),
	   .A2 (_net_7227),
	   .A1 (new_n7816_) );
   NAND4_X1 g2315 (
	   .ZN (new_n9045_),
	   .A4 (new_n7681_1_),
	   .A3 (net_7154),
	   .A2 (_net_7227),
	   .A1 (new_n7813_) );
   CLKBUF_X1 g2314 (
	   .Z (n3235),
	   .A (x1443) );
   NOR3_X1 g2313 (
	   .ZN (n3231),
	   .A3 (net_7771),
	   .A2 (new_n8911_),
	   .A1 (new_n9042_1_) );
   INV_X1 g2312 (
	   .ZN (new_n9042_1_),
	   .A (net_7770) );
   CLKBUF_X1 g2311 (
	   .Z (n3226),
	   .A (net_139) );
   OAI21_X1 g2310 (
	   .ZN (n3222),
	   .B2 (new_n6907_),
	   .B1 (new_n9039_),
	   .A (new_n9038_) );
   INV_X1 g2309 (
	   .ZN (new_n9039_),
	   .A (_net_7478) );
   NAND2_X1 g2308 (
	   .ZN (new_n9038_),
	   .A2 (new_n9037_1_),
	   .A1 (new_n6897_) );
   OAI21_X1 g2307 (
	   .ZN (new_n9037_1_),
	   .B2 (new_n9036_),
	   .B1 (new_n7034_),
	   .A (new_n9035_) );
   INV_X1 g2306 (
	   .ZN (new_n9036_),
	   .A (net_7398) );
   AOI22_X1 g2305 (
	   .ZN (new_n9035_),
	   .B2 (net_359),
	   .B1 (_net_281),
	   .A2 (_net_280),
	   .A1 (net_361) );
   NAND4_X1 g2304 (
	   .ZN (n3217),
	   .A4 (new_n9033_),
	   .A3 (new_n9027_),
	   .A2 (new_n9026_),
	   .A1 (new_n9020_) );
   AOI22_X1 g2303 (
	   .ZN (new_n9033_),
	   .B2 (_net_6110),
	   .B1 (new_n7210_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n9032_) );
   NAND4_X1 g2302 (
	   .ZN (new_n9032_),
	   .A4 (new_n9031_),
	   .A3 (new_n9030_1_),
	   .A2 (new_n9029_),
	   .A1 (new_n9028_) );
   NAND3_X1 g2301 (
	   .ZN (new_n9031_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6796) );
   NAND3_X1 g2300 (
	   .ZN (new_n9030_1_),
	   .A3 (_net_6824),
	   .A2 (net_6764),
	   .A1 (new_n7186_) );
   NAND3_X1 g2299 (
	   .ZN (new_n9029_),
	   .A3 (_net_6823),
	   .A2 (net_6732),
	   .A1 (new_n7187_) );
   NAND2_X1 g2298 (
	   .ZN (new_n9028_),
	   .A2 (net_6700),
	   .A1 (new_n7566_) );
   NAND2_X1 g2297 (
	   .ZN (new_n9027_),
	   .A2 (new_n7587_),
	   .A1 (new_n8252_) );
   NAND2_X1 g2296 (
	   .ZN (new_n9026_),
	   .A2 (new_n9025_1_),
	   .A1 (new_n7556_) );
   NAND4_X1 g2295 (
	   .ZN (new_n9025_1_),
	   .A4 (new_n9024_),
	   .A3 (new_n9023_),
	   .A2 (new_n9022_1_),
	   .A1 (new_n9021_) );
   NAND3_X1 g2294 (
	   .ZN (new_n9024_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6808) );
   NAND3_X1 g2293 (
	   .ZN (new_n9023_),
	   .A3 (_net_6824),
	   .A2 (net_6776),
	   .A1 (new_n7570_) );
   NAND3_X1 g2292 (
	   .ZN (new_n9022_1_),
	   .A3 (net_6744),
	   .A2 (_net_6823),
	   .A1 (new_n7568_) );
   NAND2_X1 g2291 (
	   .ZN (new_n9021_),
	   .A2 (net_6712),
	   .A1 (new_n7566_) );
   NAND2_X1 g2290 (
	   .ZN (new_n9020_),
	   .A2 (new_n7565_),
	   .A1 (new_n8245_1_) );
   OAI21_X1 g2289 (
	   .ZN (n3212),
	   .B2 (new_n7225_),
	   .B1 (new_n9018_),
	   .A (new_n9017_1_) );
   INV_X1 g2288 (
	   .ZN (new_n9018_),
	   .A (_net_7326) );
   NAND2_X1 g2287 (
	   .ZN (new_n9017_1_),
	   .A2 (new_n8042_1_),
	   .A1 (new_n7222_) );
   CLKBUF_X1 g2286 (
	   .Z (n3207),
	   .A (_net_7793) );
   OAI221_X1 g2285 (
	   .ZN (n3203),
	   .C2 (new_n6920_),
	   .C1 (new_n9014_1_),
	   .B2 (new_n6917_),
	   .B1 (new_n9013_),
	   .A (new_n9012_) );
   INV_X1 g2284 (
	   .ZN (new_n9014_1_),
	   .A (net_7368) );
   INV_X1 g2283 (
	   .ZN (new_n9013_),
	   .A (net_7304) );
   AOI22_X1 g2282 (
	   .ZN (new_n9012_),
	   .B2 (_net_7272),
	   .B1 (new_n6913_),
	   .A2 (net_7336),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g2281 (
	   .Z (n3199),
	   .A (net_7536) );
   AOI21_X1 g2280 (
	   .ZN (n3194),
	   .B2 (new_n7326_1_),
	   .B1 (new_n9009_),
	   .A (new_n9008_) );
   INV_X1 g2279 (
	   .ZN (new_n9009_),
	   .A (_net_7277) );
   NOR2_X1 g2278 (
	   .ZN (new_n9008_),
	   .A2 (n6376),
	   .A1 (new_n7326_1_) );
   NOR2_X1 g2277 (
	   .ZN (n6376),
	   .A2 (new_n8104_),
	   .A1 (new_n6952_1_) );
   CLKBUF_X1 g2276 (
	   .Z (n3190),
	   .A (net_6861) );
   CLKBUF_X1 g2275 (
	   .Z (n3186),
	   .A (_net_7798) );
   OAI21_X1 g2274 (
	   .ZN (n3182),
	   .B2 (new_n7111_1_),
	   .B1 (new_n7310_),
	   .A (new_n9003_) );
   NAND2_X1 g2273 (
	   .ZN (new_n9003_),
	   .A2 (new_n9002_),
	   .A1 (new_n7101_) );
   OAI221_X1 g2272 (
	   .ZN (new_n9002_),
	   .C2 (new_n7333_),
	   .C1 (new_n7105_),
	   .B2 (new_n7320_),
	   .B1 (new_n7106_),
	   .A (new_n9001_) );
   NAND2_X1 g2271 (
	   .ZN (new_n9001_),
	   .A2 (net_7238),
	   .A1 (new_n6942_) );
   CLKBUF_X1 g2270 (
	   .Z (n3178),
	   .A (net_6450) );
   CLKBUF_X1 g2269 (
	   .Z (n3174),
	   .A (_net_7815) );
   OAI21_X1 g2268 (
	   .ZN (n3170),
	   .B2 (new_n6907_),
	   .B1 (new_n8997_),
	   .A (new_n8996_) );
   INV_X1 g2267 (
	   .ZN (new_n8997_),
	   .A (_net_7470) );
   NAND2_X1 g2266 (
	   .ZN (new_n8996_),
	   .A2 (new_n7963_),
	   .A1 (new_n6897_) );
   NAND2_X1 g2265 (
	   .ZN (n3165),
	   .A2 (n4304),
	   .A1 (new_n7422_1_) );
   CLKBUF_X1 g2264 (
	   .Z (n3162),
	   .A (net_6751) );
   CLKBUF_X1 g2263 (
	   .Z (n3152),
	   .A (_net_7805) );
   OAI21_X1 g2262 (
	   .ZN (n3148),
	   .B2 (new_n7279_),
	   .B1 (new_n8991_),
	   .A (new_n8990_1_) );
   INV_X1 g2261 (
	   .ZN (new_n8991_),
	   .A (_net_7449) );
   NAND2_X1 g2260 (
	   .ZN (new_n8990_1_),
	   .A2 (new_n6904_),
	   .A1 (new_n7272_) );
   CLKBUF_X1 g2259 (
	   .Z (n3143),
	   .A (_net_7819) );
   MUX2_X1 g2258 (
	   .Z (n3139),
	   .S (new_n7609_),
	   .B (_net_7557),
	   .A (new_n7542_) );
   CLKBUF_X1 g2257 (
	   .Z (n3134),
	   .A (_net_7809) );
   OAI21_X1 g2256 (
	   .ZN (n3130),
	   .B2 (new_n7652_),
	   .B1 (new_n8985_),
	   .A (new_n8984_) );
   INV_X1 g2255 (
	   .ZN (new_n8985_),
	   .A (_net_7410) );
   NAND2_X1 g2254 (
	   .ZN (new_n8984_),
	   .A2 (new_n6935_),
	   .A1 (new_n7646_) );
   CLKBUF_X1 g2253 (
	   .Z (n3126),
	   .A (net_7387) );
   AND2_X1 g2252 (
	   .ZN (n3121),
	   .A2 (net_381),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g2251 (
	   .Z (n3117),
	   .A (_net_7824) );
   CLKBUF_X1 g2250 (
	   .Z (n3114),
	   .A (net_6743) );
   CLKBUF_X1 g2249 (
	   .Z (n3110),
	   .A (net_6473) );
   CLKBUF_X1 g2248 (
	   .Z (n3105),
	   .A (net_6396) );
   CLKBUF_X1 g2247 (
	   .Z (n3102),
	   .A (net_6706) );
   MUX2_X1 g2246 (
	   .Z (n3097),
	   .S (_net_154),
	   .B (net_324),
	   .A (_net_128) );
   AND2_X1 g2245 (
	   .ZN (n3092),
	   .A2 (_net_6280),
	   .A1 (new_n7239_) );
   NOR2_X1 g2244 (
	   .ZN (n3087),
	   .A2 (new_n8973_),
	   .A1 (new_n8972_) );
   NOR3_X1 g2243 (
	   .ZN (new_n8973_),
	   .A3 (new_n6985_),
	   .A2 (new_n7004_),
	   .A1 (new_n7013_1_) );
   NOR3_X1 g2242 (
	   .ZN (new_n8972_),
	   .A3 (new_n8218_),
	   .A2 (_net_6688),
	   .A1 (new_n7000_1_) );
   CLKBUF_X1 g2241 (
	   .Z (n3082),
	   .A (net_7799) );
   NAND2_X1 g2240 (
	   .ZN (n3078),
	   .A2 (new_n8969_),
	   .A1 (new_n8968_) );
   AOI22_X1 g2239 (
	   .ZN (new_n8969_),
	   .B2 (_net_7555),
	   .B1 (new_n6755_),
	   .A2 (_net_7619),
	   .A1 (new_n6746_1_) );
   AOI22_X1 g2238 (
	   .ZN (new_n8968_),
	   .B2 (_net_7587),
	   .B1 (new_n7350_),
	   .A2 (new_n7970_1_),
	   .A1 (_net_7651) );
   CLKBUF_X1 g2237 (
	   .Z (n3074),
	   .A (net_6717) );
   CLKBUF_X1 g2236 (
	   .Z (n3069),
	   .A (_net_7806) );
   OAI221_X1 g2235 (
	   .ZN (n3065),
	   .C2 (new_n6920_),
	   .C1 (new_n8964_),
	   .B2 (new_n6917_),
	   .B1 (new_n8963_1_),
	   .A (new_n8962_) );
   INV_X1 g2234 (
	   .ZN (new_n8964_),
	   .A (net_7374) );
   INV_X1 g2233 (
	   .ZN (new_n8963_1_),
	   .A (net_7310) );
   AOI22_X1 g2232 (
	   .ZN (new_n8962_),
	   .B2 (_net_7278),
	   .B1 (new_n6913_),
	   .A2 (net_7342),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g2231 (
	   .Z (n3061),
	   .A (net_7121) );
   NOR2_X1 g2230 (
	   .ZN (n3056),
	   .A2 (new_n8959_),
	   .A1 (new_n8958_1_) );
   XNOR2_X1 g2229 (
	   .ZN (new_n8959_),
	   .B (_net_7531),
	   .A (_net_7535) );
   NAND2_X1 g2228 (
	   .ZN (new_n8958_1_),
	   .A2 (new_n8957_),
	   .A1 (n8850) );
   XNOR2_X1 g2227 (
	   .ZN (new_n8957_),
	   .B (_net_7530),
	   .A (_net_7534) );
   XNOR2_X1 g2226 (
	   .ZN (n8850),
	   .B (_net_7533),
	   .A (net_7529) );
   CLKBUF_X1 g2225 (
	   .Z (n3052),
	   .A (net_7136) );
   MUX2_X1 g2224 (
	   .Z (n3047),
	   .S (new_n7545_),
	   .B (_net_7667),
	   .A (new_n7216_1_) );
   MUX2_X1 g2223 (
	   .Z (n3042),
	   .S (new_n7437_1_),
	   .B (_net_6023),
	   .A (_net_7823) );
   CLKBUF_X1 g2222 (
	   .Z (n3037),
	   .A (_net_7809) );
   CLKBUF_X1 g2221 (
	   .Z (n3033),
	   .A (_net_7806) );
   CLKBUF_X1 g2220 (
	   .Z (n3030),
	   .A (net_7105) );
   OAI221_X1 g2219 (
	   .ZN (n3025),
	   .C2 (new_n6920_),
	   .C1 (new_n8948_1_),
	   .B2 (new_n6917_),
	   .B1 (new_n7669_),
	   .A (new_n8947_) );
   INV_X1 g2218 (
	   .ZN (new_n8948_1_),
	   .A (_net_7363) );
   AOI22_X1 g2217 (
	   .ZN (new_n8947_),
	   .B2 (_net_7267),
	   .B1 (new_n6913_),
	   .A2 (_net_7331),
	   .A1 (new_n6911_) );
   OAI21_X1 g2216 (
	   .ZN (n3020),
	   .B2 (new_n7225_),
	   .B1 (new_n8945_),
	   .A (new_n8944_) );
   INV_X1 g2215 (
	   .ZN (new_n8945_),
	   .A (_net_7320) );
   NAND2_X1 g2214 (
	   .ZN (new_n8944_),
	   .A2 (new_n8292_),
	   .A1 (new_n7222_) );
   AND2_X1 g2213 (
	   .ZN (n3015),
	   .A2 (net_379),
	   .A1 (new_n7262_) );
   INV_X1 g2212 (
	   .ZN (n3010),
	   .A (new_n6981_) );
   NAND4_X1 g2211 (
	   .ZN (n3005),
	   .A4 (new_n8940_),
	   .A3 (new_n8934_1_),
	   .A2 (new_n8928_),
	   .A1 (new_n8927_) );
   AOI22_X1 g2210 (
	   .ZN (new_n8940_),
	   .B2 (_net_6090),
	   .B1 (new_n6985_),
	   .A2 (new_n6980_),
	   .A1 (new_n8939_1_) );
   NAND4_X1 g2209 (
	   .ZN (new_n8939_1_),
	   .A4 (new_n8938_),
	   .A3 (new_n8937_),
	   .A2 (new_n8936_),
	   .A1 (new_n8935_) );
   NAND3_X1 g2208 (
	   .ZN (new_n8938_),
	   .A3 (_net_6689),
	   .A2 (net_6661),
	   .A1 (_net_6688) );
   NAND3_X1 g2207 (
	   .ZN (new_n8937_),
	   .A3 (net_6629),
	   .A2 (_net_6689),
	   .A1 (new_n6970_) );
   NAND3_X1 g2206 (
	   .ZN (new_n8936_),
	   .A3 (net_6597),
	   .A2 (_net_6688),
	   .A1 (new_n7002_) );
   NAND2_X1 g2205 (
	   .ZN (new_n8935_),
	   .A2 (net_6565),
	   .A1 (new_n6973_) );
   NAND2_X1 g2204 (
	   .ZN (new_n8934_1_),
	   .A2 (new_n8933_),
	   .A1 (new_n7000_1_) );
   NAND4_X1 g2203 (
	   .ZN (new_n8933_),
	   .A4 (new_n8932_),
	   .A3 (new_n8931_1_),
	   .A2 (new_n8930_),
	   .A1 (new_n8929_) );
   NAND3_X1 g2202 (
	   .ZN (new_n8932_),
	   .A3 (net_6673),
	   .A2 (_net_6689),
	   .A1 (_net_6688) );
   NAND3_X1 g2201 (
	   .ZN (new_n8931_1_),
	   .A3 (_net_6689),
	   .A2 (net_6641),
	   .A1 (new_n7004_) );
   NAND3_X1 g2200 (
	   .ZN (new_n8930_),
	   .A3 (net_6609),
	   .A2 (_net_6688),
	   .A1 (new_n7002_) );
   NAND2_X1 g2199 (
	   .ZN (new_n8929_),
	   .A2 (net_6577),
	   .A1 (new_n6973_) );
   NAND2_X1 g2198 (
	   .ZN (new_n8928_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n6975_) );
   NAND2_X1 g2197 (
	   .ZN (new_n8927_),
	   .A2 (new_n7013_1_),
	   .A1 (new_n6992_) );
   OAI21_X1 g2196 (
	   .ZN (n3000),
	   .B2 (new_n8925_),
	   .B1 (new_n8920_),
	   .A (new_n8919_) );
   OAI21_X1 g2195 (
	   .ZN (new_n8925_),
	   .B2 (new_n8924_),
	   .B1 (new_n8922_1_),
	   .A (new_n8810_) );
   NOR2_X1 g2194 (
	   .ZN (new_n8924_),
	   .A2 (_net_7095),
	   .A1 (new_n8923_) );
   INV_X1 g2193 (
	   .ZN (new_n8923_),
	   .A (_net_7098) );
   NOR2_X1 g2192 (
	   .ZN (new_n8922_1_),
	   .A2 (_net_7098),
	   .A1 (new_n8921_) );
   INV_X1 g2191 (
	   .ZN (new_n8921_),
	   .A (_net_7095) );
   NAND2_X1 g2190 (
	   .ZN (new_n8920_),
	   .A2 (_net_5979),
	   .A1 (n2270) );
   INV_X1 g2189 (
	   .ZN (new_n8919_),
	   .A (_net_6038) );
   CLKBUF_X1 g2188 (
	   .Z (n2996),
	   .A (net_6438) );
   NOR3_X1 g2187 (
	   .ZN (n2991),
	   .A3 (new_n7508_),
	   .A2 (new_n8916_),
	   .A1 (new_n8915_) );
   AOI21_X1 g2186 (
	   .ZN (new_n8916_),
	   .B2 (_net_227),
	   .B1 (new_n7460_),
	   .A (_net_7531) );
   AND3_X1 g2185 (
	   .ZN (new_n8915_),
	   .A3 (_net_227),
	   .A2 (_net_7531),
	   .A1 (new_n7460_) );
   AOI21_X1 g2184 (
	   .ZN (n2986),
	   .B2 (new_n8911_),
	   .B1 (new_n8913_),
	   .A (new_n8912_1_) );
   INV_X1 g2183 (
	   .ZN (new_n8913_),
	   .A (_net_6063) );
   NOR3_X1 g2182 (
	   .ZN (new_n8912_1_),
	   .A3 (net_155),
	   .A2 (net_7767),
	   .A1 (new_n8911_) );
   INV_X1 g2181 (
	   .ZN (new_n8911_),
	   .A (_net_7791) );
   NOR2_X1 g2180 (
	   .ZN (n2981),
	   .A2 (new_n8909_),
	   .A1 (new_n8907_) );
   NOR3_X1 g2179 (
	   .ZN (new_n8909_),
	   .A3 (new_n8908_1_),
	   .A2 (_net_6553),
	   .A1 (new_n8205_) );
   NOR2_X1 g2178 (
	   .ZN (new_n8908_1_),
	   .A2 (new_n6761_1_),
	   .A1 (new_n6760_) );
   NOR3_X1 g2177 (
	   .ZN (new_n8907_),
	   .A3 (new_n6813_1_),
	   .A2 (new_n6789_),
	   .A1 (new_n6784_) );
   XNOR2_X1 g2176 (
	   .ZN (n2976),
	   .B (new_n8905_),
	   .A (new_n8410_1_) );
   NAND2_X1 g2175 (
	   .ZN (new_n8905_),
	   .A2 (net_7680),
	   .A1 (new_n7502_) );
   CLKBUF_X1 g2174 (
	   .Z (n2972),
	   .A (net_7007) );
   CLKBUF_X1 g2173 (
	   .Z (n2967),
	   .A (net_6392) );
   CLKBUF_X1 g2172 (
	   .Z (n2963),
	   .A (_net_6142) );
   NOR2_X1 g2171 (
	   .ZN (n2958),
	   .A2 (new_n8678_),
	   .A1 (new_n7035_) );
   MUX2_X1 g2170 (
	   .Z (n2953),
	   .S (new_n7609_),
	   .B (_net_7552),
	   .A (new_n8899_1_) );
   OAI21_X1 g2169 (
	   .ZN (new_n8899_1_),
	   .B2 (new_n8898_),
	   .B1 (new_n7019_),
	   .A (new_n8897_) );
   INV_X1 g2168 (
	   .ZN (new_n8898_),
	   .A (net_7536) );
   AOI22_X1 g2167 (
	   .ZN (new_n8897_),
	   .B2 (net_366),
	   .B1 (_net_292),
	   .A2 (net_368),
	   .A1 (_net_291) );
   NOR2_X1 g2166 (
	   .ZN (n2948),
	   .A2 (new_n8389_),
	   .A1 (new_n8394_) );
   CLKBUF_X1 g2165 (
	   .Z (n2944),
	   .A (net_7158) );
   CLKBUF_X1 g2164 (
	   .Z (n2939),
	   .A (_net_7816) );
   CLKBUF_X1 g2163 (
	   .Z (n2935),
	   .A (net_390) );
   AND2_X1 g2162 (
	   .ZN (n2930),
	   .A2 (_net_6220),
	   .A1 (new_n7239_) );
   CLKBUF_X1 g2161 (
	   .Z (n2926),
	   .A (net_6755) );
   CLKBUF_X1 g2160 (
	   .Z (n2922),
	   .A (net_7022) );
   NAND4_X1 g2159 (
	   .ZN (n2918),
	   .A4 (new_n8888_),
	   .A3 (new_n8887_),
	   .A2 (new_n8886_1_),
	   .A1 (new_n8884_) );
   NAND4_X1 g2158 (
	   .ZN (new_n8888_),
	   .A4 (net_7713),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   OR2_X1 g2157 (
	   .ZN (new_n8887_),
	   .A2 (new_n7339_),
	   .A1 (new_n7365_) );
   OR2_X1 g2156 (
	   .ZN (new_n8886_1_),
	   .A2 (new_n8885_),
	   .A1 (new_n7362_) );
   INV_X1 g2155 (
	   .ZN (new_n8885_),
	   .A (_net_295) );
   NOR2_X1 g2154 (
	   .ZN (new_n8884_),
	   .A2 (new_n8883_),
	   .A1 (new_n8882_1_) );
   AND2_X1 g2153 (
	   .ZN (new_n8883_),
	   .A2 (net_7742),
	   .A1 (new_n7934_) );
   NAND4_X1 g2152 (
	   .ZN (new_n8882_1_),
	   .A4 (new_n8881_),
	   .A3 (new_n8880_),
	   .A2 (new_n8879_),
	   .A1 (new_n8878_) );
   NAND4_X1 g2151 (
	   .ZN (new_n8881_),
	   .A4 (_net_178),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g2150 (
	   .ZN (new_n8880_),
	   .A3 (_net_215),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g2149 (
	   .ZN (new_n8879_),
	   .A3 (net_252),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   NAND4_X1 g2148 (
	   .ZN (new_n8878_),
	   .A4 (new_n7354_1_),
	   .A3 (net_152),
	   .A2 (x1261),
	   .A1 (new_n7370_) );
   NOR2_X1 g2147 (
	   .ZN (n2913),
	   .A2 (new_n7494_),
	   .A1 (new_n6952_1_) );
   CLKBUF_X1 g2146 (
	   .Z (n2908),
	   .A (_net_7814) );
   NOR2_X1 g2145 (
	   .ZN (n2904),
	   .A2 (new_n6900_),
	   .A1 (new_n8543_) );
   AOI21_X1 g2144 (
	   .ZN (n2900),
	   .B2 (new_n8873_1_),
	   .B1 (new_n8872_),
	   .A (new_n7428_) );
   INV_X1 g2143 (
	   .ZN (new_n8873_1_),
	   .A (_net_7722) );
   INV_X1 g2142 (
	   .ZN (new_n8872_),
	   .A (net_5992) );
   CLKBUF_X1 g2141 (
	   .Z (n2895),
	   .A (_net_5972) );
   MUX2_X1 g2140 (
	   .Z (n2890),
	   .S (new_n7609_),
	   .B (_net_7572),
	   .A (n615) );
   CLKBUF_X1 g2139 (
	   .Z (n2885),
	   .A (_net_7816) );
   CLKBUF_X1 g2138 (
	   .Z (n2882),
	   .A (net_7547) );
   CLKBUF_X1 g2137 (
	   .Z (n2877),
	   .A (_net_6068) );
   CLKBUF_X1 g2136 (
	   .Z (n2873),
	   .A (net_6578) );
   CLKBUF_X1 g2135 (
	   .Z (n2869),
	   .A (net_6478) );
   CLKBUF_X1 g2134 (
	   .Z (n2864),
	   .A (_net_6070) );
   CLKBUF_X1 g2133 (
	   .Z (n2860),
	   .A (net_7236) );
   OAI21_X1 g2132 (
	   .ZN (n2855),
	   .B2 (new_n7736_),
	   .B1 (new_n8861_),
	   .A (new_n8860_1_) );
   INV_X1 g2131 (
	   .ZN (new_n8861_),
	   .A (_net_7501) );
   NAND2_X1 g2130 (
	   .ZN (new_n8860_1_),
	   .A2 (new_n8859_),
	   .A1 (new_n7733_) );
   OAI21_X1 g2129 (
	   .ZN (new_n8859_),
	   .B2 (new_n8858_),
	   .B1 (new_n7034_),
	   .A (new_n8857_) );
   INV_X1 g2128 (
	   .ZN (new_n8858_),
	   .A (net_7389) );
   AOI22_X1 g2127 (
	   .ZN (new_n8857_),
	   .B2 (net_350),
	   .B1 (_net_281),
	   .A2 (_net_280),
	   .A1 (net_352) );
   AND2_X1 g2126 (
	   .ZN (n2850),
	   .A2 (net_376),
	   .A1 (new_n7262_) );
   OAI21_X1 g2125 (
	   .ZN (n2845),
	   .B2 (new_n6957_1_),
	   .B1 (new_n8854_),
	   .A (new_n8853_) );
   INV_X1 g2124 (
	   .ZN (new_n8854_),
	   .A (_net_7261) );
   NAND2_X1 g2123 (
	   .ZN (new_n8853_),
	   .A2 (new_n8852_),
	   .A1 (new_n6949_) );
   OAI221_X1 g2122 (
	   .ZN (new_n8852_),
	   .C2 (new_n7105_),
	   .C1 (new_n8103_),
	   .B2 (new_n7106_),
	   .B1 (new_n7104_),
	   .A (new_n8851_) );
   NAND2_X1 g2121 (
	   .ZN (new_n8851_),
	   .A2 (net_7245),
	   .A1 (new_n6942_) );
   CLKBUF_X1 g2120 (
	   .Z (n2840),
	   .A (_net_7801) );
   OAI21_X1 g2119 (
	   .ZN (n2836),
	   .B2 (new_n6823_),
	   .B1 (new_n8091_),
	   .A (new_n8848_) );
   NAND2_X1 g2118 (
	   .ZN (new_n8848_),
	   .A2 (_net_6029),
	   .A1 (new_n6823_) );
   NAND3_X1 g2117 (
	   .ZN (n2831),
	   .A3 (new_n8846_),
	   .A2 (new_n8840_1_),
	   .A1 (new_n8831_1_) );
   AOI22_X1 g2116 (
	   .ZN (new_n8846_),
	   .B2 (new_n8180_),
	   .B1 (net_7084),
	   .A2 (new_n8845_1_),
	   .A1 (new_n7060_) );
   NAND4_X1 g2115 (
	   .ZN (new_n8845_1_),
	   .A4 (new_n8844_),
	   .A3 (new_n8843_),
	   .A2 (new_n8842_),
	   .A1 (new_n8841_) );
   NAND3_X1 g2114 (
	   .ZN (new_n8844_),
	   .A3 (net_7068),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   NAND3_X1 g2113 (
	   .ZN (new_n8843_),
	   .A3 (net_7036),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g2112 (
	   .ZN (new_n8842_),
	   .A3 (_net_7093),
	   .A2 (net_7004),
	   .A1 (new_n7075_) );
   NAND2_X1 g2111 (
	   .ZN (new_n8841_),
	   .A2 (net_6972),
	   .A1 (new_n7063_) );
   AND3_X1 g2110 (
	   .ZN (new_n8840_1_),
	   .A3 (new_n8839_),
	   .A2 (new_n8838_),
	   .A1 (new_n8832_) );
   NAND2_X1 g2109 (
	   .ZN (new_n8839_),
	   .A2 (_net_6156),
	   .A1 (new_n7092_) );
   NAND2_X1 g2108 (
	   .ZN (new_n8838_),
	   .A2 (new_n7070_),
	   .A1 (new_n8837_) );
   NAND4_X1 g2107 (
	   .ZN (new_n8837_),
	   .A4 (new_n8836_),
	   .A3 (new_n8835_1_),
	   .A2 (new_n8834_),
	   .A1 (new_n8833_) );
   NAND3_X1 g2106 (
	   .ZN (new_n8836_),
	   .A3 (_net_7093),
	   .A2 (net_7070),
	   .A1 (_net_7094) );
   NAND3_X1 g2105 (
	   .ZN (new_n8835_1_),
	   .A3 (net_7038),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g2104 (
	   .ZN (new_n8834_),
	   .A3 (net_7006),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   NAND2_X1 g2103 (
	   .ZN (new_n8833_),
	   .A2 (net_6974),
	   .A1 (new_n7063_) );
   NAND2_X1 g2102 (
	   .ZN (new_n8832_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n8670_) );
   AND3_X1 g2101 (
	   .ZN (new_n8831_1_),
	   .A3 (new_n8830_),
	   .A2 (new_n8829_),
	   .A1 (new_n8828_) );
   NAND4_X1 g2100 (
	   .ZN (new_n8830_),
	   .A4 (new_n7044_),
	   .A3 (_net_7092),
	   .A2 (net_7052),
	   .A1 (new_n8158_) );
   NAND4_X1 g2099 (
	   .ZN (new_n8829_),
	   .A4 (new_n7052_),
	   .A3 (net_6988),
	   .A2 (_net_7092),
	   .A1 (new_n8158_) );
   NAND4_X1 g2098 (
	   .ZN (new_n8828_),
	   .A4 (new_n7050_),
	   .A3 (net_7020),
	   .A2 (_net_7092),
	   .A1 (new_n8155_) );
   CLKBUF_X1 g2097 (
	   .Z (n2827),
	   .A (net_7153) );
   CLKBUF_X1 g2096 (
	   .Z (n2823),
	   .A (net_7024) );
   CLKBUF_X1 g2095 (
	   .Z (n2819),
	   .A (net_6579) );
   CLKBUF_X1 g2094 (
	   .Z (n2814),
	   .A (_net_7812) );
   NAND2_X1 g2093 (
	   .ZN (n2810),
	   .A2 (new_n8822_),
	   .A1 (new_n8821_) );
   AOI22_X1 g2092 (
	   .ZN (new_n8822_),
	   .B2 (net_7518),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7486) );
   AOI22_X1 g2091 (
	   .ZN (new_n8821_),
	   .B2 (_net_7422),
	   .B1 (new_n7298_),
	   .A2 (net_7454),
	   .A1 (new_n7296_) );
   CLKBUF_X1 g2090 (
	   .Z (n2805),
	   .A (x1374) );
   CLKBUF_X1 g2089 (
	   .Z (n2801),
	   .A (_net_7797) );
   NAND2_X1 g2088 (
	   .ZN (n2797),
	   .A2 (new_n8817_),
	   .A1 (new_n8816_) );
   AOI22_X1 g2087 (
	   .ZN (new_n8817_),
	   .B2 (_net_7554),
	   .B1 (new_n6755_),
	   .A2 (_net_7618),
	   .A1 (new_n6746_1_) );
   AOI22_X1 g2086 (
	   .ZN (new_n8816_),
	   .B2 (_net_7586),
	   .B1 (new_n7350_),
	   .A2 (new_n7970_1_),
	   .A1 (_net_7650) );
   CLKBUF_X1 g2085 (
	   .Z (n2792),
	   .A (net_7802) );
   CLKBUF_X1 g2084 (
	   .Z (n2788),
	   .A (_net_7801) );
   AND2_X1 g2083 (
	   .ZN (n2784),
	   .A2 (net_343),
	   .A1 (new_n7102_1_) );
   CLKBUF_X1 g2082 (
	   .Z (n2781),
	   .A (net_6880) );
   XNOR2_X1 g2081 (
	   .ZN (n2776),
	   .B (new_n8438_1_),
	   .A (new_n8810_) );
   XNOR2_X1 g2080 (
	   .ZN (new_n8810_),
	   .B (_net_7097),
	   .A (_net_7094) );
   MUX2_X1 g2079 (
	   .Z (n2771),
	   .S (new_n7437_1_),
	   .B (_net_6022),
	   .A (_net_7822) );
   CLKBUF_X1 g2078 (
	   .Z (n2767),
	   .A (net_7108) );
   CLKBUF_X1 g2077 (
	   .Z (n2762),
	   .A (_net_7823) );
   NAND3_X1 g2076 (
	   .ZN (n2758),
	   .A3 (new_n8805_1_),
	   .A2 (new_n8804_),
	   .A1 (new_n8795_) );
   AOI22_X1 g2075 (
	   .ZN (new_n8805_1_),
	   .B2 (new_n7136_),
	   .B1 (net_6680),
	   .A2 (new_n7916_1_),
	   .A1 (new_n7013_1_) );
   AND3_X1 g2074 (
	   .ZN (new_n8804_),
	   .A3 (new_n8803_),
	   .A2 (new_n8802_),
	   .A1 (new_n8801_) );
   NAND2_X1 g2073 (
	   .ZN (new_n8803_),
	   .A2 (_net_6097),
	   .A1 (new_n6985_) );
   NAND2_X1 g2072 (
	   .ZN (new_n8802_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n7910_) );
   NAND2_X1 g2071 (
	   .ZN (new_n8801_),
	   .A2 (new_n6980_),
	   .A1 (new_n8800_1_) );
   NAND4_X1 g2070 (
	   .ZN (new_n8800_1_),
	   .A4 (new_n8799_),
	   .A3 (new_n8798_),
	   .A2 (new_n8797_1_),
	   .A1 (new_n8796_) );
   NAND3_X1 g2069 (
	   .ZN (new_n8799_),
	   .A3 (_net_6689),
	   .A2 (net_6668),
	   .A1 (_net_6688) );
   NAND3_X1 g2068 (
	   .ZN (new_n8798_),
	   .A3 (_net_6689),
	   .A2 (net_6636),
	   .A1 (new_n7004_) );
   NAND3_X1 g2067 (
	   .ZN (new_n8797_1_),
	   .A3 (net_6604),
	   .A2 (_net_6688),
	   .A1 (new_n7002_) );
   NAND2_X1 g2066 (
	   .ZN (new_n8796_),
	   .A2 (net_6572),
	   .A1 (new_n6973_) );
   AND3_X1 g2065 (
	   .ZN (new_n8795_),
	   .A3 (new_n8794_),
	   .A2 (new_n8793_1_),
	   .A1 (new_n8792_) );
   NAND4_X1 g2064 (
	   .ZN (new_n8794_),
	   .A4 (new_n6987_),
	   .A3 (net_6648),
	   .A2 (_net_6687),
	   .A1 (new_n7118_) );
   NAND4_X1 g2063 (
	   .ZN (new_n8793_1_),
	   .A4 (new_n6990_1_),
	   .A3 (_net_6687),
	   .A2 (net_6584),
	   .A1 (new_n7115_) );
   NAND4_X1 g2062 (
	   .ZN (new_n8792_),
	   .A4 (new_n6989_),
	   .A3 (_net_6687),
	   .A2 (net_6616),
	   .A1 (new_n7115_) );
   OAI221_X1 g2061 (
	   .ZN (n2753),
	   .C2 (new_n7312_1_),
	   .C1 (new_n8790_),
	   .B2 (new_n7986_),
	   .B1 (new_n8789_),
	   .A (new_n8788_1_) );
   INV_X1 g2060 (
	   .ZN (new_n8790_),
	   .A (_net_7289) );
   INV_X1 g2059 (
	   .ZN (new_n8789_),
	   .A (_net_7353) );
   AOI22_X1 g2058 (
	   .ZN (new_n8788_1_),
	   .B2 (_net_7257),
	   .B1 (new_n6913_),
	   .A2 (_net_7321),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g2057 (
	   .Z (n2748),
	   .A (_net_7823) );
   CLKBUF_X1 g2056 (
	   .Z (n2745),
	   .A (net_6725) );
   CLKBUF_X1 g2055 (
	   .Z (n2741),
	   .A (net_6586) );
   CLKBUF_X1 g2054 (
	   .Z (n2737),
	   .A (net_7708) );
   OAI21_X1 g2053 (
	   .ZN (n2732),
	   .B2 (new_n7225_),
	   .B1 (new_n8782_),
	   .A (new_n8781_) );
   INV_X1 g2052 (
	   .ZN (new_n8782_),
	   .A (_net_7314) );
   NAND2_X1 g2051 (
	   .ZN (new_n8781_),
	   .A2 (new_n8780_1_),
	   .A1 (new_n7222_) );
   OAI21_X1 g2050 (
	   .ZN (new_n8780_1_),
	   .B2 (new_n8779_),
	   .B1 (new_n6951_),
	   .A (new_n8778_) );
   INV_X1 g2049 (
	   .ZN (new_n8779_),
	   .A (net_7234) );
   AOI22_X1 g2048 (
	   .ZN (new_n8778_),
	   .B2 (net_328),
	   .B1 (_net_269),
	   .A2 (_net_270),
	   .A1 (net_326) );
   CLKBUF_X1 g2047 (
	   .Z (n2727),
	   .A (net_6381) );
   MUX2_X1 g2046 (
	   .Z (n2723),
	   .S (new_n7538_),
	   .B (_net_280),
	   .A (_net_7803) );
   NAND2_X1 g2045 (
	   .ZN (n2718),
	   .A2 (new_n8774_),
	   .A1 (new_n8773_) );
   AOI22_X1 g2044 (
	   .ZN (new_n8774_),
	   .B2 (new_n6751_),
	   .B1 (_net_7560),
	   .A2 (_net_7656),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g2043 (
	   .ZN (new_n8773_),
	   .B2 (_net_7592),
	   .B1 (new_n7350_),
	   .A2 (new_n6746_1_),
	   .A1 (_net_7624) );
   MUX2_X1 g2042 (
	   .Z (n2713),
	   .S (_net_154),
	   .B (net_322),
	   .A (_net_126) );
   CLKBUF_X1 g2041 (
	   .Z (n2709),
	   .A (net_6969) );
   CLKBUF_X1 g2040 (
	   .Z (n2705),
	   .A (net_6434) );
   CLKBUF_X1 g2039 (
	   .Z (n2701),
	   .A (net_6981) );
   NAND2_X1 g2038 (
	   .ZN (n2696),
	   .A2 (new_n8767_1_),
	   .A1 (new_n8766_) );
   INV_X1 g2037 (
	   .ZN (new_n8767_1_),
	   .A (new_n7565_) );
   OAI21_X1 g2036 (
	   .ZN (new_n8766_),
	   .B2 (new_n7210_),
	   .B1 (new_n8765_),
	   .A (_net_6822) );
   NOR2_X1 g2035 (
	   .ZN (new_n8765_),
	   .A2 (new_n7200_),
	   .A1 (new_n8764_) );
   INV_X1 g2034 (
	   .ZN (new_n8764_),
	   .A (new_n7553_1_) );
   CLKBUF_X1 g2033 (
	   .Z (n2692),
	   .A (net_7393) );
   AND2_X1 g2032 (
	   .ZN (n2687),
	   .A2 (new_n8761_),
	   .A1 (new_n8760_) );
   INV_X1 g2031 (
	   .ZN (new_n8761_),
	   .A (x906) );
   AOI211_X1 g2030 (
	   .ZN (new_n8760_),
	   .C2 (new_n8759_),
	   .C1 (new_n8758_),
	   .B (new_n8754_),
	   .A (new_n8753_1_) );
   AOI21_X1 g2029 (
	   .ZN (new_n8759_),
	   .B2 (new_n8757_1_),
	   .B1 (new_n8756_),
	   .A (_net_5980) );
   OAI21_X1 g2028 (
	   .ZN (new_n8758_),
	   .B2 (new_n8757_1_),
	   .B1 (new_n8756_),
	   .A (new_n8755_) );
   INV_X1 g2027 (
	   .ZN (new_n8757_1_),
	   .A (_net_5982) );
   NOR2_X1 g2026 (
	   .ZN (new_n8756_),
	   .A2 (_net_6043),
	   .A1 (_net_5981) );
   INV_X1 g2025 (
	   .ZN (new_n8755_),
	   .A (_net_6044) );
   INV_X1 g2024 (
	   .ZN (new_n8754_),
	   .A (_net_6039) );
   INV_X1 g2023 (
	   .ZN (new_n8753_1_),
	   .A (_net_6045) );
   CLKBUF_X1 g2022 (
	   .Z (n2682),
	   .A (_net_7822) );
   CLKBUF_X1 g2021 (
	   .Z (n2679),
	   .A (net_6964) );
   CLKBUF_X1 g2020 (
	   .Z (n2675),
	   .A (net_6890) );
   CLKBUF_X1 g2019 (
	   .Z (n2670),
	   .A (_net_6134) );
   NAND2_X1 g2018 (
	   .ZN (n2665),
	   .A2 (new_n8747_),
	   .A1 (new_n8727_) );
   AND4_X1 g2017 (
	   .ZN (new_n8747_),
	   .A4 (new_n8746_),
	   .A3 (new_n8745_),
	   .A2 (new_n8739_1_),
	   .A1 (new_n8733_) );
   NAND2_X1 g2016 (
	   .ZN (new_n8746_),
	   .A2 (_net_6121),
	   .A1 (new_n7210_) );
   NAND2_X1 g2015 (
	   .ZN (new_n8745_),
	   .A2 (new_n7587_),
	   .A1 (new_n8744_) );
   NAND4_X1 g2014 (
	   .ZN (new_n8744_),
	   .A4 (new_n8743_1_),
	   .A3 (new_n8742_),
	   .A2 (new_n8741_),
	   .A1 (new_n8740_) );
   NAND3_X1 g2013 (
	   .ZN (new_n8743_1_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6805) );
   NAND3_X1 g2012 (
	   .ZN (new_n8742_),
	   .A3 (_net_6824),
	   .A2 (net_6773),
	   .A1 (new_n7570_) );
   NAND3_X1 g2011 (
	   .ZN (new_n8741_),
	   .A3 (_net_6823),
	   .A2 (net_6741),
	   .A1 (new_n7568_) );
   NAND2_X1 g2010 (
	   .ZN (new_n8740_),
	   .A2 (net_6709),
	   .A1 (new_n7566_) );
   NAND2_X1 g2009 (
	   .ZN (new_n8739_1_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n8738_) );
   NAND4_X1 g2008 (
	   .ZN (new_n8738_),
	   .A4 (new_n8737_),
	   .A3 (new_n8736_),
	   .A2 (new_n8735_),
	   .A1 (new_n8734_1_) );
   NAND3_X1 g2007 (
	   .ZN (new_n8737_),
	   .A3 (net_6807),
	   .A2 (_net_6824),
	   .A1 (_net_6823) );
   NAND3_X1 g2006 (
	   .ZN (new_n8736_),
	   .A3 (net_6775),
	   .A2 (_net_6824),
	   .A1 (new_n7570_) );
   NAND3_X1 g2005 (
	   .ZN (new_n8735_),
	   .A3 (_net_6823),
	   .A2 (net_6743),
	   .A1 (new_n7568_) );
   NAND2_X1 g2004 (
	   .ZN (new_n8734_1_),
	   .A2 (net_6711),
	   .A1 (new_n7566_) );
   NAND2_X1 g2003 (
	   .ZN (new_n8733_),
	   .A2 (new_n8732_),
	   .A1 (new_n7565_) );
   NAND4_X1 g2002 (
	   .ZN (new_n8732_),
	   .A4 (new_n8731_),
	   .A3 (new_n8730_1_),
	   .A2 (new_n8729_),
	   .A1 (new_n8728_) );
   NAND3_X1 g2001 (
	   .ZN (new_n8731_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6803) );
   NAND3_X1 g2000 (
	   .ZN (new_n8730_1_),
	   .A3 (_net_6824),
	   .A2 (net_6771),
	   .A1 (new_n7570_) );
   NAND3_X1 g1999 (
	   .ZN (new_n8729_),
	   .A3 (_net_6823),
	   .A2 (net_6739),
	   .A1 (new_n7568_) );
   NAND2_X1 g1998 (
	   .ZN (new_n8728_),
	   .A2 (net_6707),
	   .A1 (new_n7566_) );
   AND4_X1 g1997 (
	   .ZN (new_n8727_),
	   .A4 (new_n8726_),
	   .A3 (new_n8725_1_),
	   .A2 (new_n8724_),
	   .A1 (new_n8723_) );
   NAND4_X1 g1996 (
	   .ZN (new_n8726_),
	   .A4 (new_n7194_1_),
	   .A3 (net_6755),
	   .A2 (_net_6822),
	   .A1 (new_n7559_) );
   NAND4_X1 g1995 (
	   .ZN (new_n8725_1_),
	   .A4 (new_n7191_),
	   .A3 (net_6787),
	   .A2 (_net_6822),
	   .A1 (new_n7560_) );
   NAND3_X1 g1994 (
	   .ZN (new_n8724_),
	   .A3 (new_n7189_),
	   .A2 (net_6819),
	   .A1 (new_n7555_) );
   NAND3_X1 g1993 (
	   .ZN (new_n8723_),
	   .A3 (new_n7196_),
	   .A2 (net_6723),
	   .A1 (new_n7556_) );
   CLKBUF_X1 g1992 (
	   .Z (n2660),
	   .A (net_149) );
   CLKBUF_X1 g1991 (
	   .Z (n2656),
	   .A (net_6606) );
   OAI221_X1 g1990 (
	   .ZN (n2651),
	   .C2 (new_n7312_1_),
	   .C1 (new_n8719_),
	   .B2 (new_n7986_),
	   .B1 (new_n8718_),
	   .A (new_n8717_) );
   INV_X1 g1989 (
	   .ZN (new_n8719_),
	   .A (net_7313) );
   INV_X1 g1988 (
	   .ZN (new_n8718_),
	   .A (net_7377) );
   AOI22_X1 g1987 (
	   .ZN (new_n8717_),
	   .B2 (_net_7281),
	   .B1 (new_n6913_),
	   .A2 (net_7345),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g1986 (
	   .Z (n2647),
	   .A (net_6588) );
   CLKBUF_X1 g1985 (
	   .Z (n2642),
	   .A (_net_6145) );
   NAND2_X1 g1984 (
	   .ZN (n2637),
	   .A2 (new_n8713_),
	   .A1 (new_n8712_) );
   AOI22_X1 g1983 (
	   .ZN (new_n8713_),
	   .B2 (_net_7579),
	   .B1 (new_n6755_),
	   .A2 (net_7611),
	   .A1 (new_n6743_) );
   AOI22_X1 g1982 (
	   .ZN (new_n8712_),
	   .B2 (net_7643),
	   .B1 (new_n8009_),
	   .A2 (new_n7970_1_),
	   .A1 (net_7675) );
   AND2_X1 g1981 (
	   .ZN (n2632),
	   .A2 (_net_5924),
	   .A1 (net_5858) );
   CLKBUF_X1 g1980 (
	   .Z (n2627),
	   .A (_net_6126) );
   CLKBUF_X1 g1979 (
	   .Z (n2622),
	   .A (_net_7822) );
   CLKBUF_X1 g1978 (
	   .Z (n2618),
	   .A (_net_7793) );
   CLKBUF_X1 g1977 (
	   .Z (n2615),
	   .A (net_6967) );
   CLKBUF_X1 g1976 (
	   .Z (n2610),
	   .A (_net_6181) );
   CLKBUF_X1 g1975 (
	   .Z (n2605),
	   .A (_net_7818) );
   CLKBUF_X1 g1974 (
	   .Z (n2601),
	   .A (_net_7822) );
   CLKBUF_X1 g1973 (
	   .Z (n2597),
	   .A (_net_7797) );
   CLKBUF_X1 g1972 (
	   .Z (n2594),
	   .A (net_6390) );
   NOR2_X1 g1971 (
	   .ZN (n2590),
	   .A2 (new_n7090_),
	   .A1 (new_n8700_) );
   INV_X1 g1970 (
	   .ZN (new_n8700_),
	   .A (_net_5979) );
   NOR2_X1 g1969 (
	   .ZN (n2585),
	   .A2 (x868),
	   .A1 (new_n8698_1_) );
   NAND2_X1 g1968 (
	   .ZN (new_n8698_1_),
	   .A2 (_net_284),
	   .A1 (n3827) );
   OAI221_X1 g1967 (
	   .ZN (n2580),
	   .C2 (new_n7303_),
	   .C1 (new_n8696_),
	   .B2 (new_n7306_),
	   .B1 (new_n8566_),
	   .A (new_n8695_) );
   INV_X1 g1966 (
	   .ZN (new_n8696_),
	   .A (_net_7479) );
   AOI22_X1 g1965 (
	   .ZN (new_n8695_),
	   .B2 (_net_7415),
	   .B1 (new_n7298_),
	   .A2 (_net_7447),
	   .A1 (new_n8694_1_) );
   BUF_X4 g1964 (
	   .Z (new_n8694_1_),
	   .A (new_n7295_) );
   OAI221_X1 g1963 (
	   .ZN (n2575),
	   .C2 (new_n7312_1_),
	   .C1 (new_n8692_),
	   .B2 (new_n7986_),
	   .B1 (new_n8691_),
	   .A (new_n8690_) );
   INV_X1 g1962 (
	   .ZN (new_n8692_),
	   .A (net_7302) );
   INV_X1 g1961 (
	   .ZN (new_n8691_),
	   .A (net_7366) );
   AOI22_X1 g1960 (
	   .ZN (new_n8690_),
	   .B2 (_net_7270),
	   .B1 (new_n6913_),
	   .A2 (net_7334),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g1959 (
	   .Z (n2570),
	   .A (_net_7798) );
   MUX2_X1 g1958 (
	   .Z (n2566),
	   .S (new_n7545_),
	   .B (_net_7663),
	   .A (new_n8687_) );
   OAI21_X1 g1957 (
	   .ZN (new_n8687_),
	   .B2 (new_n8686_),
	   .B1 (new_n7019_),
	   .A (new_n8685_1_) );
   INV_X1 g1956 (
	   .ZN (new_n8686_),
	   .A (net_7551) );
   AOI22_X1 g1955 (
	   .ZN (new_n8685_1_),
	   .B2 (_net_291),
	   .B1 (net_383),
	   .A2 (_net_292),
	   .A1 (net_381) );
   CLKBUF_X1 g1954 (
	   .Z (n2561),
	   .A (net_6390) );
   CLKBUF_X1 g1953 (
	   .Z (n2556),
	   .A (_net_7819) );
   OAI21_X1 g1952 (
	   .ZN (n2552),
	   .B2 (new_n7279_),
	   .B1 (new_n8681_1_),
	   .A (new_n8680_) );
   INV_X1 g1951 (
	   .ZN (new_n8681_1_),
	   .A (_net_7445) );
   NAND2_X1 g1950 (
	   .ZN (new_n8680_),
	   .A2 (new_n8679_),
	   .A1 (new_n7272_) );
   OAI221_X1 g1949 (
	   .ZN (new_n8679_),
	   .C2 (new_n8678_),
	   .C1 (new_n6901_),
	   .B2 (new_n6902_1_),
	   .B1 (new_n7594_),
	   .A (new_n8677_) );
   INV_X1 g1948 (
	   .ZN (new_n8678_),
	   .A (net_358) );
   NAND2_X1 g1947 (
	   .ZN (new_n8677_),
	   .A2 (net_7397),
	   .A1 (new_n6889_) );
   NOR2_X1 g1946 (
	   .ZN (n2547),
	   .A2 (new_n7104_),
	   .A1 (new_n8675_) );
   BUF_X4 g1945 (
	   .Z (new_n8675_),
	   .A (new_n6952_1_) );
   CLKBUF_X1 g1944 (
	   .Z (n2543),
	   .A (net_7807) );
   CLKBUF_X1 g1943 (
	   .Z (n2539),
	   .A (_net_7797) );
   NAND3_X1 g1942 (
	   .ZN (n2534),
	   .A3 (new_n8671_1_),
	   .A2 (new_n8665_),
	   .A1 (new_n8651_) );
   AOI22_X1 g1941 (
	   .ZN (new_n8671_1_),
	   .B2 (new_n8180_),
	   .B1 (net_7088),
	   .A2 (new_n8670_),
	   .A1 (new_n7060_) );
   NAND4_X1 g1940 (
	   .ZN (new_n8670_),
	   .A4 (new_n8669_),
	   .A3 (new_n8668_),
	   .A2 (new_n8667_),
	   .A1 (new_n8666_1_) );
   NAND3_X1 g1939 (
	   .ZN (new_n8669_),
	   .A3 (net_7072),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   NAND3_X1 g1938 (
	   .ZN (new_n8668_),
	   .A3 (net_7040),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g1937 (
	   .ZN (new_n8667_),
	   .A3 (net_7008),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   NAND2_X1 g1936 (
	   .ZN (new_n8666_1_),
	   .A2 (net_6976),
	   .A1 (new_n7063_) );
   AND3_X1 g1935 (
	   .ZN (new_n8665_),
	   .A3 (new_n8664_),
	   .A2 (new_n8663_),
	   .A1 (new_n8657_) );
   NAND2_X1 g1934 (
	   .ZN (new_n8664_),
	   .A2 (_net_6160),
	   .A1 (new_n7092_) );
   NAND2_X1 g1933 (
	   .ZN (new_n8663_),
	   .A2 (new_n7070_),
	   .A1 (new_n8662_1_) );
   NAND4_X1 g1932 (
	   .ZN (new_n8662_1_),
	   .A4 (new_n8661_),
	   .A3 (new_n8660_),
	   .A2 (new_n8659_),
	   .A1 (new_n8658_1_) );
   NAND3_X1 g1931 (
	   .ZN (new_n8661_),
	   .A3 (net_7074),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   NAND3_X1 g1930 (
	   .ZN (new_n8660_),
	   .A3 (net_7042),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g1929 (
	   .ZN (new_n8659_),
	   .A3 (_net_7093),
	   .A2 (net_7010),
	   .A1 (new_n7075_) );
   NAND2_X1 g1928 (
	   .ZN (new_n8658_1_),
	   .A2 (net_6978),
	   .A1 (new_n7063_) );
   NAND2_X1 g1927 (
	   .ZN (new_n8657_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n8656_) );
   NAND4_X1 g1926 (
	   .ZN (new_n8656_),
	   .A4 (new_n8655_),
	   .A3 (new_n8654_1_),
	   .A2 (new_n8653_),
	   .A1 (new_n8652_) );
   NAND3_X1 g1925 (
	   .ZN (new_n8655_),
	   .A3 (net_7076),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   NAND3_X1 g1924 (
	   .ZN (new_n8654_1_),
	   .A3 (net_7044),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g1923 (
	   .ZN (new_n8653_),
	   .A3 (net_7012),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   NAND2_X1 g1922 (
	   .ZN (new_n8652_),
	   .A2 (net_6980),
	   .A1 (new_n7063_) );
   AND3_X1 g1921 (
	   .ZN (new_n8651_),
	   .A3 (new_n8650_1_),
	   .A2 (new_n8649_),
	   .A1 (new_n8648_) );
   NAND4_X1 g1920 (
	   .ZN (new_n8650_1_),
	   .A4 (new_n7044_),
	   .A3 (net_7056),
	   .A2 (_net_7092),
	   .A1 (new_n8158_) );
   NAND4_X1 g1919 (
	   .ZN (new_n8649_),
	   .A4 (new_n7052_),
	   .A3 (net_6992),
	   .A2 (_net_7092),
	   .A1 (new_n8155_) );
   NAND4_X1 g1918 (
	   .ZN (new_n8648_),
	   .A4 (new_n7050_),
	   .A3 (_net_7092),
	   .A2 (net_7024),
	   .A1 (new_n8155_) );
   OAI21_X1 g1917 (
	   .ZN (n2529),
	   .B2 (new_n7652_),
	   .B1 (new_n8646_),
	   .A (new_n8645_1_) );
   INV_X1 g1916 (
	   .ZN (new_n8646_),
	   .A (_net_7419) );
   NAND2_X1 g1915 (
	   .ZN (new_n8645_1_),
	   .A2 (new_n8280_1_),
	   .A1 (new_n7646_) );
   OAI221_X1 g1914 (
	   .ZN (n2524),
	   .C2 (new_n7312_1_),
	   .C1 (new_n8643_),
	   .B2 (new_n7986_),
	   .B1 (new_n8642_),
	   .A (new_n8641_1_) );
   INV_X1 g1913 (
	   .ZN (new_n8643_),
	   .A (net_7305) );
   INV_X1 g1912 (
	   .ZN (new_n8642_),
	   .A (net_7369) );
   AOI22_X1 g1911 (
	   .ZN (new_n8641_1_),
	   .B2 (_net_7273),
	   .B1 (new_n6913_),
	   .A2 (net_7337),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g1910 (
	   .Z (n2519),
	   .A (_net_7795) );
   AOI21_X1 g1909 (
	   .ZN (n2515),
	   .B2 (new_n7344_1_),
	   .B1 (new_n7343_),
	   .A (new_n7208_) );
   NAND2_X1 g1908 (
	   .ZN (n2510),
	   .A2 (new_n8637_1_),
	   .A1 (new_n8636_) );
   AOI22_X1 g1907 (
	   .ZN (new_n8637_1_),
	   .B2 (_net_7574),
	   .B1 (new_n6755_),
	   .A2 (net_7606),
	   .A1 (new_n6743_) );
   AOI22_X1 g1906 (
	   .ZN (new_n8636_),
	   .B2 (net_7638),
	   .B1 (new_n8009_),
	   .A2 (new_n7970_1_),
	   .A1 (net_7670) );
   MUX2_X1 g1905 (
	   .Z (n2505),
	   .S (new_n7285_),
	   .B (_net_7704),
	   .A (_net_7806) );
   AND2_X1 g1904 (
	   .ZN (n2500),
	   .A2 (net_377),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g1903 (
	   .Z (n2496),
	   .A (_net_7805) );
   CLKBUF_X1 g1902 (
	   .Z (n2493),
	   .A (net_6435) );
   CLKBUF_X1 g1901 (
	   .Z (n2488),
	   .A (net_7799) );
   NAND2_X1 g1900 (
	   .ZN (n2484),
	   .A2 (new_n8629_),
	   .A1 (new_n8628_1_) );
   AOI22_X1 g1899 (
	   .ZN (new_n8629_),
	   .B2 (net_7528),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7496) );
   AOI22_X1 g1898 (
	   .ZN (new_n8628_1_),
	   .B2 (_net_7432),
	   .B1 (new_n7298_),
	   .A2 (net_7464),
	   .A1 (new_n7296_) );
   OAI21_X1 g1897 (
	   .ZN (n2479),
	   .B2 (new_n7258_),
	   .B1 (new_n8626_),
	   .A (new_n8625_1_) );
   INV_X1 g1896 (
	   .ZN (new_n8626_),
	   .A (_net_7294) );
   NAND2_X1 g1895 (
	   .ZN (new_n8625_1_),
	   .A2 (new_n8042_1_),
	   .A1 (new_n7252_1_) );
   CLKBUF_X1 g1894 (
	   .Z (n2474),
	   .A (_net_7810) );
   NAND2_X1 g1893 (
	   .ZN (n2470),
	   .A2 (new_n8622_),
	   .A1 (new_n8612_1_) );
   AND4_X1 g1892 (
	   .ZN (new_n8622_),
	   .A4 (new_n8621_1_),
	   .A3 (new_n8620_),
	   .A2 (new_n8619_),
	   .A1 (new_n8618_) );
   NAND2_X1 g1891 (
	   .ZN (new_n8621_1_),
	   .A2 (_net_6118),
	   .A1 (new_n7210_) );
   NAND2_X1 g1890 (
	   .ZN (new_n8620_),
	   .A2 (new_n7587_),
	   .A1 (new_n7573_) );
   NAND2_X1 g1889 (
	   .ZN (new_n8619_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n7585_) );
   NAND2_X1 g1888 (
	   .ZN (new_n8618_),
	   .A2 (new_n8617_),
	   .A1 (new_n7565_) );
   NAND4_X1 g1887 (
	   .ZN (new_n8617_),
	   .A4 (new_n8616_1_),
	   .A3 (new_n8615_),
	   .A2 (new_n8614_),
	   .A1 (new_n8613_) );
   NAND3_X1 g1886 (
	   .ZN (new_n8616_1_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6800) );
   NAND3_X1 g1885 (
	   .ZN (new_n8615_),
	   .A3 (_net_6824),
	   .A2 (net_6768),
	   .A1 (new_n7570_) );
   NAND3_X1 g1884 (
	   .ZN (new_n8614_),
	   .A3 (_net_6823),
	   .A2 (net_6736),
	   .A1 (new_n7568_) );
   NAND2_X1 g1883 (
	   .ZN (new_n8613_),
	   .A2 (net_6704),
	   .A1 (new_n7566_) );
   AND4_X1 g1882 (
	   .ZN (new_n8612_1_),
	   .A4 (new_n8611_),
	   .A3 (new_n8610_),
	   .A2 (new_n8609_),
	   .A1 (new_n8608_) );
   NAND4_X1 g1881 (
	   .ZN (new_n8611_),
	   .A4 (new_n7194_1_),
	   .A3 (net_6752),
	   .A2 (_net_6822),
	   .A1 (new_n7560_) );
   NAND4_X1 g1880 (
	   .ZN (new_n8610_),
	   .A4 (new_n7191_),
	   .A3 (_net_6822),
	   .A2 (net_6784),
	   .A1 (new_n7560_) );
   NAND3_X1 g1879 (
	   .ZN (new_n8609_),
	   .A3 (new_n7189_),
	   .A2 (net_6816),
	   .A1 (new_n7555_) );
   NAND3_X1 g1878 (
	   .ZN (new_n8608_),
	   .A3 (new_n7196_),
	   .A2 (net_6720),
	   .A1 (new_n7556_) );
   CLKBUF_X1 g1877 (
	   .Z (n2465),
	   .A (_net_7818) );
   CLKBUF_X1 g1876 (
	   .Z (n2462),
	   .A (net_6426) );
   MUX2_X1 g1875 (
	   .Z (n2457),
	   .S (new_n7437_1_),
	   .B (_net_5984),
	   .A (_net_7793) );
   CLKBUF_X1 g1874 (
	   .Z (n2452),
	   .A (_net_7824) );
   CLKBUF_X1 g1873 (
	   .Z (n2448),
	   .A (net_6392) );
   NOR2_X1 g1872 (
	   .ZN (n2444),
	   .A2 (new_n8601_),
	   .A1 (new_n8599_) );
   XNOR2_X1 g1871 (
	   .ZN (new_n8601_),
	   .B (new_n8600_),
	   .A (new_n8402_) );
   INV_X1 g1870 (
	   .ZN (new_n8600_),
	   .A (_net_6963) );
   NAND4_X1 g1869 (
	   .ZN (new_n8599_),
	   .A4 (new_n8598_1_),
	   .A3 (new_n8597_),
	   .A2 (new_n8596_),
	   .A1 (new_n8594_) );
   NAND2_X1 g1868 (
	   .ZN (new_n8598_1_),
	   .A2 (_net_6962),
	   .A1 (new_n8593_1_) );
   OR2_X1 g1867 (
	   .ZN (new_n8597_),
	   .A2 (_net_6957),
	   .A1 (n9778) );
   OAI21_X1 g1866 (
	   .ZN (new_n8596_),
	   .B2 (new_n6827_),
	   .B1 (n9778),
	   .A (_net_6957) );
   XNOR2_X1 g1865 (
	   .ZN (n9778),
	   .B (_net_6958),
	   .A (net_6961) );
   OR2_X1 g1864 (
	   .ZN (new_n8594_),
	   .A2 (_net_6962),
	   .A1 (new_n8593_1_) );
   NAND2_X1 g1863 (
	   .ZN (new_n8593_1_),
	   .A2 (new_n6880_),
	   .A1 (new_n8592_) );
   OAI21_X1 g1862 (
	   .ZN (new_n8592_),
	   .B2 (new_n6848_),
	   .B1 (new_n8591_),
	   .A (new_n6846_) );
   INV_X1 g1861 (
	   .ZN (new_n8591_),
	   .A (_net_6957) );
   CLKBUF_X1 g1860 (
	   .Z (n2440),
	   .A (net_7240) );
   MUX2_X1 g1859 (
	   .Z (n2435),
	   .S (new_n7538_),
	   .B (_net_279),
	   .A (net_7802) );
   AOI21_X1 g1858 (
	   .ZN (n2430),
	   .B2 (new_n7739_),
	   .B1 (new_n8587_),
	   .A (new_n8586_) );
   INV_X1 g1857 (
	   .ZN (new_n8587_),
	   .A (_net_7431) );
   NOR2_X1 g1856 (
	   .ZN (new_n8586_),
	   .A2 (n1752),
	   .A1 (new_n7739_) );
   CLKBUF_X1 g1855 (
	   .Z (n2426),
	   .A (net_6833) );
   CLKBUF_X1 g1854 (
	   .Z (n2422),
	   .A (net_7016) );
   CLKBUF_X1 g1853 (
	   .Z (n2417),
	   .A (_net_7818) );
   NAND3_X1 g1852 (
	   .ZN (n2414),
	   .A3 (new_n8581_),
	   .A2 (new_n8580_),
	   .A1 (new_n8572_) );
   NAND4_X1 g1851 (
	   .ZN (new_n8581_),
	   .A4 (_net_7695),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR3_X1 g1850 (
	   .ZN (new_n8580_),
	   .A3 (new_n8579_),
	   .A2 (new_n8575_1_),
	   .A1 (new_n8573_) );
   NAND3_X1 g1849 (
	   .ZN (new_n8579_),
	   .A3 (new_n8578_1_),
	   .A2 (new_n8577_),
	   .A1 (new_n8576_) );
   NAND4_X1 g1848 (
	   .ZN (new_n8578_1_),
	   .A4 (net_160),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g1847 (
	   .ZN (new_n8577_),
	   .A3 (net_197),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g1846 (
	   .ZN (new_n8576_),
	   .A3 (net_234),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   OAI22_X1 g1845 (
	   .ZN (new_n8575_1_),
	   .B2 (new_n7378_),
	   .B1 (new_n8415_1_),
	   .A2 (new_n8574_),
	   .A1 (new_n7374_) );
   INV_X1 g1844 (
	   .ZN (new_n8574_),
	   .A (_net_118) );
   AND4_X1 g1843 (
	   .ZN (new_n8573_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7369_),
	   .A1 (_net_6032) );
   NOR2_X1 g1842 (
	   .ZN (new_n8572_),
	   .A2 (new_n8571_),
	   .A1 (new_n8569_) );
   NOR2_X1 g1841 (
	   .ZN (new_n8571_),
	   .A2 (new_n8570_1_),
	   .A1 (new_n7366_) );
   INV_X1 g1840 (
	   .ZN (new_n8570_1_),
	   .A (_net_5988) );
   NOR2_X1 g1839 (
	   .ZN (new_n8569_),
	   .A2 (new_n8568_),
	   .A1 (new_n7362_) );
   INV_X1 g1838 (
	   .ZN (new_n8568_),
	   .A (_net_271) );
   OAI21_X1 g1837 (
	   .ZN (n2409),
	   .B2 (new_n7736_),
	   .B1 (new_n8566_),
	   .A (new_n8565_1_) );
   INV_X1 g1836 (
	   .ZN (new_n8566_),
	   .A (_net_7511) );
   NAND2_X1 g1835 (
	   .ZN (new_n8565_1_),
	   .A2 (new_n7595_),
	   .A1 (new_n7733_) );
   AND2_X1 g1834 (
	   .ZN (n2404),
	   .A2 (net_378),
	   .A1 (new_n7262_) );
   CLKBUF_X1 g1833 (
	   .Z (n2399),
	   .A (_net_7793) );
   OAI221_X1 g1832 (
	   .ZN (n2395),
	   .C2 (new_n6920_),
	   .C1 (new_n8561_1_),
	   .B2 (new_n6917_),
	   .B1 (new_n8560_),
	   .A (new_n8559_) );
   INV_X1 g1831 (
	   .ZN (new_n8561_1_),
	   .A (net_7373) );
   INV_X1 g1830 (
	   .ZN (new_n8560_),
	   .A (net_7309) );
   AOI22_X1 g1829 (
	   .ZN (new_n8559_),
	   .B2 (_net_7277),
	   .B1 (new_n6913_),
	   .A2 (net_7341),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g1828 (
	   .Z (n2391),
	   .A (net_6576) );
   NAND4_X1 g1827 (
	   .ZN (n2386),
	   .A4 (new_n8556_),
	   .A3 (new_n8555_),
	   .A2 (new_n8554_),
	   .A1 (new_n8548_) );
   NAND2_X1 g1826 (
	   .ZN (new_n8556_),
	   .A2 (new_n7837_),
	   .A1 (new_n7698_) );
   NAND2_X1 g1825 (
	   .ZN (new_n8555_),
	   .A2 (new_n7701_),
	   .A1 (new_n7685_) );
   NAND2_X1 g1824 (
	   .ZN (new_n8554_),
	   .A2 (new_n8553_),
	   .A1 (new_n8026_) );
   NAND4_X1 g1823 (
	   .ZN (new_n8553_),
	   .A4 (new_n8552_1_),
	   .A3 (new_n8551_),
	   .A2 (new_n8550_),
	   .A1 (new_n8549_1_) );
   NAND3_X1 g1822 (
	   .ZN (new_n8552_1_),
	   .A3 (net_7212),
	   .A2 (_net_7228),
	   .A1 (_net_7229) );
   NAND3_X1 g1821 (
	   .ZN (new_n8551_),
	   .A3 (net_7180),
	   .A2 (_net_7229),
	   .A1 (new_n7823_) );
   NAND3_X1 g1820 (
	   .ZN (new_n8550_),
	   .A3 (_net_7228),
	   .A2 (net_7148),
	   .A1 (new_n7821_) );
   NAND2_X1 g1819 (
	   .ZN (new_n8549_1_),
	   .A2 (net_7116),
	   .A1 (new_n7819_) );
   AOI22_X1 g1818 (
	   .ZN (new_n8548_),
	   .B2 (new_n7694_),
	   .B1 (_net_6169),
	   .A2 (new_n7690_),
	   .A1 (new_n8547_) );
   NAND2_X1 g1817 (
	   .ZN (new_n8547_),
	   .A2 (new_n8546_),
	   .A1 (new_n8545_) );
   AOI22_X1 g1816 (
	   .ZN (new_n8546_),
	   .B2 (net_7104),
	   .B1 (new_n7819_),
	   .A2 (net_7136),
	   .A1 (new_n7680_) );
   AOI22_X1 g1815 (
	   .ZN (new_n8545_),
	   .B2 (net_7168),
	   .B1 (new_n7677_),
	   .A2 (new_n7676_1_),
	   .A1 (net_7200) );
   NOR2_X1 g1814 (
	   .ZN (n2381),
	   .A2 (new_n6903_),
	   .A1 (new_n8543_) );
   BUF_X4 g1813 (
	   .Z (new_n8543_),
	   .A (new_n7035_) );
   AOI21_X1 g1812 (
	   .ZN (n2377),
	   .B2 (new_n8541_),
	   .B1 (new_n8540_1_),
	   .A (new_n7428_) );
   INV_X1 g1811 (
	   .ZN (new_n8541_),
	   .A (_net_154) );
   INV_X1 g1810 (
	   .ZN (new_n8540_1_),
	   .A (_net_7720) );
   CLKBUF_X1 g1809 (
	   .Z (n2373),
	   .A (net_6397) );
   CLKBUF_X1 g1808 (
	   .Z (n2370),
	   .A (net_6593) );
   NAND3_X1 g1807 (
	   .ZN (n2365),
	   .A3 (new_n8536_),
	   .A2 (new_n8530_),
	   .A1 (new_n8516_) );
   AOI22_X1 g1806 (
	   .ZN (new_n8536_),
	   .B2 (new_n8180_),
	   .B1 (net_7091),
	   .A2 (new_n8535_1_),
	   .A1 (new_n7060_) );
   NAND4_X1 g1805 (
	   .ZN (new_n8535_1_),
	   .A4 (new_n8534_),
	   .A3 (new_n8533_),
	   .A2 (new_n8532_),
	   .A1 (new_n8531_1_) );
   NAND3_X1 g1804 (
	   .ZN (new_n8534_),
	   .A3 (net_7075),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   NAND3_X1 g1803 (
	   .ZN (new_n8533_),
	   .A3 (net_7043),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g1802 (
	   .ZN (new_n8532_),
	   .A3 (net_7011),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   NAND2_X1 g1801 (
	   .ZN (new_n8531_1_),
	   .A2 (net_6979),
	   .A1 (new_n7063_) );
   AND3_X1 g1800 (
	   .ZN (new_n8530_),
	   .A3 (new_n8529_),
	   .A2 (new_n8528_),
	   .A1 (new_n8522_1_) );
   NAND2_X1 g1799 (
	   .ZN (new_n8529_),
	   .A2 (_net_6163),
	   .A1 (new_n7092_) );
   NAND2_X1 g1798 (
	   .ZN (new_n8528_),
	   .A2 (new_n7088_),
	   .A1 (new_n8527_) );
   NAND4_X1 g1797 (
	   .ZN (new_n8527_),
	   .A4 (new_n8526_1_),
	   .A3 (new_n8525_),
	   .A2 (new_n8524_),
	   .A1 (new_n8523_) );
   NAND3_X1 g1796 (
	   .ZN (new_n8526_1_),
	   .A3 (net_7079),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   NAND3_X1 g1795 (
	   .ZN (new_n8525_),
	   .A3 (net_7047),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g1794 (
	   .ZN (new_n8524_),
	   .A3 (net_7015),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   NAND2_X1 g1793 (
	   .ZN (new_n8523_),
	   .A2 (net_6983),
	   .A1 (new_n7063_) );
   NAND2_X1 g1792 (
	   .ZN (new_n8522_1_),
	   .A2 (new_n7070_),
	   .A1 (new_n8521_) );
   NAND4_X1 g1791 (
	   .ZN (new_n8521_),
	   .A4 (new_n8520_),
	   .A3 (new_n8519_),
	   .A2 (new_n8518_),
	   .A1 (new_n8517_1_) );
   NAND3_X1 g1790 (
	   .ZN (new_n8520_),
	   .A3 (net_7077),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   NAND3_X1 g1789 (
	   .ZN (new_n8519_),
	   .A3 (net_7045),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g1788 (
	   .ZN (new_n8518_),
	   .A3 (net_7013),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   NAND2_X1 g1787 (
	   .ZN (new_n8517_1_),
	   .A2 (net_6981),
	   .A1 (new_n7063_) );
   AND3_X1 g1786 (
	   .ZN (new_n8516_),
	   .A3 (new_n8515_),
	   .A2 (new_n8514_),
	   .A1 (new_n8513_1_) );
   NAND4_X1 g1785 (
	   .ZN (new_n8515_),
	   .A4 (new_n7044_),
	   .A3 (net_7059),
	   .A2 (_net_7092),
	   .A1 (new_n8158_) );
   NAND4_X1 g1784 (
	   .ZN (new_n8514_),
	   .A4 (new_n7052_),
	   .A3 (_net_7092),
	   .A2 (net_6995),
	   .A1 (new_n8155_) );
   NAND4_X1 g1783 (
	   .ZN (new_n8513_1_),
	   .A4 (new_n7050_),
	   .A3 (net_7027),
	   .A2 (_net_7092),
	   .A1 (new_n8155_) );
   CLKBUF_X1 g1782 (
	   .Z (n2360),
	   .A (_net_7812) );
   CLKBUF_X1 g1781 (
	   .Z (n2355),
	   .A (_net_6101) );
   CLKBUF_X1 g1780 (
	   .Z (n2350),
	   .A (net_142) );
   CLKBUF_X1 g1779 (
	   .Z (n2347),
	   .A (net_6849) );
   CLKBUF_X1 g1778 (
	   .Z (n2342),
	   .A (_net_7806) );
   CLKBUF_X1 g1777 (
	   .Z (n2338),
	   .A (_net_7820) );
   AOI21_X1 g1776 (
	   .ZN (n2334),
	   .B2 (new_n8505_),
	   .B1 (new_n6959_),
	   .A (new_n7428_) );
   INV_X1 g1775 (
	   .ZN (new_n8505_),
	   .A (_net_7747) );
   NAND3_X1 g1774 (
	   .ZN (n2329),
	   .A3 (new_n8503_),
	   .A2 (new_n8497_),
	   .A1 (new_n8483_) );
   AOI22_X1 g1773 (
	   .ZN (new_n8503_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6947),
	   .A2 (new_n8502_),
	   .A1 (new_n6879_) );
   NAND4_X1 g1772 (
	   .ZN (new_n8502_),
	   .A4 (new_n8501_),
	   .A3 (new_n8500_),
	   .A2 (new_n8499_1_),
	   .A1 (new_n8498_) );
   NAND3_X1 g1771 (
	   .ZN (new_n8501_),
	   .A3 (_net_6958),
	   .A2 (_net_6959),
	   .A1 (net_6931) );
   NAND3_X1 g1770 (
	   .ZN (new_n8500_),
	   .A3 (_net_6959),
	   .A2 (net_6899),
	   .A1 (new_n6831_1_) );
   NAND3_X1 g1769 (
	   .ZN (new_n8499_1_),
	   .A3 (_net_6958),
	   .A2 (net_6867),
	   .A1 (new_n6846_) );
   NAND2_X1 g1768 (
	   .ZN (new_n8498_),
	   .A2 (net_6835),
	   .A1 (new_n6844_) );
   AND3_X1 g1767 (
	   .ZN (new_n8497_),
	   .A3 (new_n8496_),
	   .A2 (new_n8495_),
	   .A1 (new_n8489_) );
   NAND2_X1 g1766 (
	   .ZN (new_n8496_),
	   .A2 (_net_6134),
	   .A1 (new_n6869_) );
   NAND2_X1 g1765 (
	   .ZN (new_n8495_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n8494_1_) );
   NAND4_X1 g1764 (
	   .ZN (new_n8494_1_),
	   .A4 (new_n8493_),
	   .A3 (new_n8492_),
	   .A2 (new_n8491_1_),
	   .A1 (new_n8490_) );
   NAND3_X1 g1763 (
	   .ZN (new_n8493_),
	   .A3 (_net_6958),
	   .A2 (_net_6959),
	   .A1 (net_6933) );
   NAND3_X1 g1762 (
	   .ZN (new_n8492_),
	   .A3 (_net_6959),
	   .A2 (net_6901),
	   .A1 (new_n6848_) );
   NAND3_X1 g1761 (
	   .ZN (new_n8491_1_),
	   .A3 (_net_6958),
	   .A2 (net_6869),
	   .A1 (new_n6846_) );
   NAND2_X1 g1760 (
	   .ZN (new_n8490_),
	   .A2 (net_6837),
	   .A1 (new_n6844_) );
   NAND2_X1 g1759 (
	   .ZN (new_n8489_),
	   .A2 (new_n6854_),
	   .A1 (new_n8488_) );
   NAND4_X1 g1758 (
	   .ZN (new_n8488_),
	   .A4 (new_n8487_),
	   .A3 (new_n8486_1_),
	   .A2 (new_n8485_),
	   .A1 (new_n8484_) );
   NAND3_X1 g1757 (
	   .ZN (new_n8487_),
	   .A3 (_net_6958),
	   .A2 (_net_6959),
	   .A1 (net_6935) );
   NAND3_X1 g1756 (
	   .ZN (new_n8486_1_),
	   .A3 (_net_6959),
	   .A2 (net_6903),
	   .A1 (new_n6848_) );
   NAND3_X1 g1755 (
	   .ZN (new_n8485_),
	   .A3 (net_6871),
	   .A2 (_net_6958),
	   .A1 (new_n6846_) );
   NAND2_X1 g1754 (
	   .ZN (new_n8484_),
	   .A2 (net_6839),
	   .A1 (new_n6844_) );
   AND3_X1 g1753 (
	   .ZN (new_n8483_),
	   .A3 (new_n8482_),
	   .A2 (new_n8481_1_),
	   .A1 (new_n8480_) );
   NAND4_X1 g1752 (
	   .ZN (new_n8482_),
	   .A4 (new_n6841_),
	   .A3 (_net_6957),
	   .A2 (net_6915),
	   .A1 (new_n6838_) );
   NAND4_X1 g1751 (
	   .ZN (new_n8481_1_),
	   .A4 (new_n6836_1_),
	   .A3 (net_6851),
	   .A2 (_net_6957),
	   .A1 (new_n6838_) );
   NAND4_X1 g1750 (
	   .ZN (new_n8480_),
	   .A4 (new_n6833_),
	   .A3 (_net_6957),
	   .A2 (net_6883),
	   .A1 (new_n6830_) );
   CLKBUF_X1 g1749 (
	   .Z (n2324),
	   .A (net_6398) );
   CLKBUF_X1 g1748 (
	   .Z (n2321),
	   .A (net_7159) );
   CLKBUF_X1 g1747 (
	   .Z (n2316),
	   .A (_net_7800) );
   MUX2_X1 g1746 (
	   .Z (n2312),
	   .S (new_n7609_),
	   .B (_net_7556),
	   .A (new_n8475_) );
   OAI21_X1 g1745 (
	   .ZN (new_n8475_),
	   .B2 (new_n8474_),
	   .B1 (new_n7019_),
	   .A (new_n8473_) );
   INV_X1 g1744 (
	   .ZN (new_n8474_),
	   .A (net_7540) );
   AOI22_X1 g1743 (
	   .ZN (new_n8473_),
	   .B2 (_net_292),
	   .B1 (net_370),
	   .A2 (_net_291),
	   .A1 (net_372) );
   CLKBUF_X1 g1742 (
	   .Z (n2307),
	   .A (_net_7824) );
   AND2_X1 g1741 (
	   .ZN (n2303),
	   .A2 (_net_6186),
	   .A1 (new_n7239_) );
   NAND2_X1 g1740 (
	   .ZN (n2298),
	   .A2 (new_n8469_),
	   .A1 (new_n8468_) );
   INV_X1 g1739 (
	   .ZN (new_n8469_),
	   .A (_net_6015) );
   NAND2_X1 g1738 (
	   .ZN (new_n8468_),
	   .A2 (_net_5968),
	   .A1 (new_n7207_1_) );
   CLKBUF_X1 g1737 (
	   .Z (n2293),
	   .A (_net_6170) );
   CLKBUF_X1 g1736 (
	   .Z (n2288),
	   .A (_net_7805) );
   CLKBUF_X1 g1735 (
	   .Z (n2284),
	   .A (net_6397) );
   AOI21_X1 g1734 (
	   .ZN (n2280),
	   .B2 (new_n8463_),
	   .B1 (new_n7766_),
	   .A (new_n7428_) );
   INV_X1 g1733 (
	   .ZN (new_n8463_),
	   .A (_net_7748) );
   NAND3_X1 g1732 (
	   .ZN (n2275),
	   .A3 (new_n8461_),
	   .A2 (new_n8460_),
	   .A1 (new_n8446_) );
   AOI22_X1 g1731 (
	   .ZN (new_n8461_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6952),
	   .A2 (new_n7716_),
	   .A1 (new_n6879_) );
   AND3_X1 g1730 (
	   .ZN (new_n8460_),
	   .A3 (new_n8459_1_),
	   .A2 (new_n8458_),
	   .A1 (new_n8452_) );
   NAND2_X1 g1729 (
	   .ZN (new_n8459_1_),
	   .A2 (_net_6139),
	   .A1 (new_n6869_) );
   NAND2_X1 g1728 (
	   .ZN (new_n8458_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n8457_) );
   NAND4_X1 g1727 (
	   .ZN (new_n8457_),
	   .A4 (new_n8456_),
	   .A3 (new_n8455_1_),
	   .A2 (new_n8454_),
	   .A1 (new_n8453_) );
   NAND3_X1 g1726 (
	   .ZN (new_n8456_),
	   .A3 (_net_6958),
	   .A2 (_net_6959),
	   .A1 (net_6938) );
   NAND3_X1 g1725 (
	   .ZN (new_n8455_1_),
	   .A3 (_net_6959),
	   .A2 (net_6906),
	   .A1 (new_n6848_) );
   NAND3_X1 g1724 (
	   .ZN (new_n8454_),
	   .A3 (_net_6958),
	   .A2 (net_6874),
	   .A1 (new_n6846_) );
   NAND2_X1 g1723 (
	   .ZN (new_n8453_),
	   .A2 (net_6842),
	   .A1 (new_n6844_) );
   NAND2_X1 g1722 (
	   .ZN (new_n8452_),
	   .A2 (new_n6854_),
	   .A1 (new_n8451_1_) );
   NAND4_X1 g1721 (
	   .ZN (new_n8451_1_),
	   .A4 (new_n8450_),
	   .A3 (new_n8449_),
	   .A2 (new_n8448_),
	   .A1 (new_n8447_1_) );
   NAND3_X1 g1720 (
	   .ZN (new_n8450_),
	   .A3 (_net_6958),
	   .A2 (_net_6959),
	   .A1 (net_6940) );
   NAND3_X1 g1719 (
	   .ZN (new_n8449_),
	   .A3 (net_6908),
	   .A2 (_net_6959),
	   .A1 (new_n6848_) );
   NAND3_X1 g1718 (
	   .ZN (new_n8448_),
	   .A3 (net_6876),
	   .A2 (_net_6958),
	   .A1 (new_n6846_) );
   NAND2_X1 g1717 (
	   .ZN (new_n8447_1_),
	   .A2 (net_6844),
	   .A1 (new_n6844_) );
   AND3_X1 g1716 (
	   .ZN (new_n8446_),
	   .A3 (new_n8445_),
	   .A2 (new_n8444_),
	   .A1 (new_n8443_1_) );
   NAND4_X1 g1715 (
	   .ZN (new_n8445_),
	   .A4 (new_n6841_),
	   .A3 (_net_6957),
	   .A2 (net_6920),
	   .A1 (new_n6838_) );
   NAND4_X1 g1714 (
	   .ZN (new_n8444_),
	   .A4 (new_n6836_1_),
	   .A3 (_net_6957),
	   .A2 (net_6856),
	   .A1 (new_n6830_) );
   NAND4_X1 g1713 (
	   .ZN (new_n8443_1_),
	   .A4 (new_n6833_),
	   .A3 (_net_6957),
	   .A2 (net_6888),
	   .A1 (new_n6830_) );
   INV_X1 g1712 (
	   .ZN (n2270),
	   .A (new_n8441_) );
   NAND2_X1 g1711 (
	   .ZN (new_n8441_),
	   .A2 (new_n8440_),
	   .A1 (new_n8438_1_) );
   NAND2_X1 g1710 (
	   .ZN (new_n8440_),
	   .A2 (_net_7093),
	   .A1 (new_n8439_) );
   INV_X1 g1709 (
	   .ZN (new_n8439_),
	   .A (net_7096) );
   NAND2_X1 g1708 (
	   .ZN (new_n8438_1_),
	   .A2 (net_7096),
	   .A1 (new_n7077_1_) );
   OAI21_X1 g1707 (
	   .ZN (n2265),
	   .B2 (new_n7652_),
	   .B1 (new_n8436_),
	   .A (new_n8435_1_) );
   INV_X1 g1706 (
	   .ZN (new_n8436_),
	   .A (_net_7401) );
   NAND2_X1 g1705 (
	   .ZN (new_n8435_1_),
	   .A2 (new_n7874_),
	   .A1 (new_n7646_) );
   AND2_X1 g1704 (
	   .ZN (n2260),
	   .A2 (net_377),
	   .A1 (new_n7747_) );
   XOR2_X1 g1703 (
	   .Z (n2251),
	   .B (_net_6402),
	   .A (net_6403) );
   NAND3_X1 g1702 (
	   .ZN (n2247),
	   .A3 (new_n8431_),
	   .A2 (new_n8430_1_),
	   .A1 (new_n8421_) );
   NAND4_X1 g1701 (
	   .ZN (new_n8431_),
	   .A4 (_net_7704),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR3_X1 g1700 (
	   .ZN (new_n8430_1_),
	   .A3 (new_n8429_),
	   .A2 (new_n8425_),
	   .A1 (new_n8422_1_) );
   NAND3_X1 g1699 (
	   .ZN (new_n8429_),
	   .A3 (new_n8428_),
	   .A2 (new_n8427_),
	   .A1 (new_n8426_1_) );
   NAND4_X1 g1698 (
	   .ZN (new_n8428_),
	   .A4 (net_169),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g1697 (
	   .ZN (new_n8427_),
	   .A3 (net_206),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g1696 (
	   .ZN (new_n8426_1_),
	   .A3 (net_243),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   OAI22_X1 g1695 (
	   .ZN (new_n8425_),
	   .B2 (new_n7378_),
	   .B1 (new_n8424_),
	   .A2 (new_n8423_),
	   .A1 (new_n7374_) );
   INV_X1 g1694 (
	   .ZN (new_n8424_),
	   .A (_net_7733) );
   INV_X1 g1693 (
	   .ZN (new_n8423_),
	   .A (_net_127) );
   AND4_X1 g1692 (
	   .ZN (new_n8422_1_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7369_),
	   .A1 (_net_6044) );
   NOR2_X1 g1691 (
	   .ZN (new_n8421_),
	   .A2 (new_n8420_),
	   .A1 (new_n8418_1_) );
   NOR2_X1 g1690 (
	   .ZN (new_n8420_),
	   .A2 (new_n8419_),
	   .A1 (new_n7366_) );
   INV_X1 g1689 (
	   .ZN (new_n8419_),
	   .A (_net_6000) );
   NOR2_X1 g1688 (
	   .ZN (new_n8418_1_),
	   .A2 (new_n7509_1_),
	   .A1 (new_n7362_) );
   AOI21_X1 g1687 (
	   .ZN (n2242),
	   .B2 (new_n8416_),
	   .B1 (new_n8415_1_),
	   .A (new_n7428_) );
   INV_X1 g1686 (
	   .ZN (new_n8416_),
	   .A (_net_5994) );
   INV_X1 g1685 (
	   .ZN (new_n8415_1_),
	   .A (_net_7724) );
   NOR3_X1 g1684 (
	   .ZN (n2237),
	   .A3 (x1231),
	   .A2 (x1215),
	   .A1 (new_n7182_1_) );
   NOR2_X1 g1683 (
	   .ZN (n2232),
	   .A2 (new_n8412_),
	   .A1 (new_n8411_) );
   XNOR2_X1 g1682 (
	   .ZN (new_n8412_),
	   .B (_net_7682),
	   .A (_net_7686) );
   NAND2_X1 g1681 (
	   .ZN (new_n8411_),
	   .A2 (new_n8410_1_),
	   .A1 (n4405) );
   XNOR2_X1 g1680 (
	   .ZN (new_n8410_1_),
	   .B (_net_7685),
	   .A (_net_7681) );
   XNOR2_X1 g1679 (
	   .ZN (n4405),
	   .B (net_7680),
	   .A (_net_7684) );
   NAND2_X1 g1678 (
	   .ZN (n2227),
	   .A2 (new_n8407_),
	   .A1 (new_n8403_) );
   NAND3_X1 g1677 (
	   .ZN (new_n8407_),
	   .A3 (new_n8406_),
	   .A2 (new_n8405_1_),
	   .A1 (new_n8404_) );
   NAND2_X1 g1676 (
	   .ZN (new_n8406_),
	   .A2 (new_n8400_),
	   .A1 (new_n6872_1_) );
   INV_X1 g1675 (
	   .ZN (new_n8405_1_),
	   .A (new_n8401_1_) );
   NOR2_X1 g1674 (
	   .ZN (new_n8404_),
	   .A2 (new_n6827_),
	   .A1 (new_n6826_1_) );
   AOI22_X1 g1673 (
	   .ZN (new_n8403_),
	   .B2 (_net_6960),
	   .B1 (new_n6869_),
	   .A2 (new_n6830_),
	   .A1 (new_n8402_) );
   AOI22_X1 g1672 (
	   .ZN (new_n8402_),
	   .B2 (new_n6880_),
	   .B1 (new_n8400_),
	   .A2 (_net_6957),
	   .A1 (new_n8401_1_) );
   NOR2_X1 g1671 (
	   .ZN (new_n8401_1_),
	   .A2 (new_n8400_),
	   .A1 (new_n6872_1_) );
   INV_X1 g1670 (
	   .ZN (new_n8400_),
	   .A (_net_6960) );
   AND2_X1 g1669 (
	   .ZN (n2222),
	   .A2 (_net_5984),
	   .A1 (_net_5963) );
   CLKBUF_X1 g1668 (
	   .Z (n2218),
	   .A (net_6456) );
   OAI21_X1 g1667 (
	   .ZN (n2213),
	   .B2 (new_n8396_1_),
	   .B1 (new_n8392_1_),
	   .A (new_n7744_) );
   NAND2_X1 g1666 (
	   .ZN (new_n8396_1_),
	   .A2 (new_n8395_),
	   .A1 (new_n8393_) );
   INV_X1 g1665 (
	   .ZN (new_n8395_),
	   .A (new_n8394_) );
   NOR2_X1 g1664 (
	   .ZN (new_n8394_),
	   .A2 (_net_6823),
	   .A1 (new_n8304_) );
   XNOR2_X1 g1663 (
	   .ZN (new_n8393_),
	   .B (_net_6824),
	   .A (_net_6827) );
   OR4_X1 g1662 (
	   .ZN (new_n8392_1_),
	   .A4 (new_n8391_),
	   .A3 (new_n8390_),
	   .A2 (new_n8389_),
	   .A1 (new_n8305_) );
   NOR2_X1 g1661 (
	   .ZN (new_n8391_),
	   .A2 (_net_6828),
	   .A1 (_net_6825) );
   AND2_X1 g1660 (
	   .ZN (new_n8390_),
	   .A2 (_net_6828),
	   .A1 (_net_6825) );
   NOR2_X1 g1659 (
	   .ZN (new_n8389_),
	   .A2 (net_6826),
	   .A1 (new_n7570_) );
   NOR2_X1 g1658 (
	   .ZN (n2208),
	   .A2 (new_n8387_1_),
	   .A1 (new_n8386_) );
   INV_X1 g1657 (
	   .ZN (new_n8387_1_),
	   .A (new_n7364_) );
   NAND3_X1 g1656 (
	   .ZN (new_n8386_),
	   .A3 (new_n7395_1_),
	   .A2 (x1231),
	   .A1 (new_n7183_) );
   CLKBUF_X1 g1655 (
	   .Z (n2203),
	   .A (_net_7796) );
   OAI221_X1 g1654 (
	   .ZN (n2199),
	   .C2 (new_n8383_),
	   .C1 (new_n8024_1_),
	   .B2 (new_n7692_),
	   .B1 (new_n7821_),
	   .A (new_n8380_) );
   NAND2_X1 g1653 (
	   .ZN (new_n8383_),
	   .A2 (new_n7843_),
	   .A1 (new_n8382_1_) );
   NAND2_X1 g1652 (
	   .ZN (new_n8382_1_),
	   .A2 (new_n7821_),
	   .A1 (new_n8381_) );
   NAND2_X1 g1651 (
	   .ZN (new_n8381_),
	   .A2 (_net_7228),
	   .A1 (_net_7227) );
   OAI21_X1 g1650 (
	   .ZN (new_n8380_),
	   .B2 (new_n7678_),
	   .B1 (new_n7681_1_),
	   .A (new_n8379_) );
   NOR2_X1 g1649 (
	   .ZN (new_n8379_),
	   .A2 (new_n7810_1_),
	   .A1 (new_n7687_) );
   NAND3_X1 g1648 (
	   .ZN (n2194),
	   .A3 (new_n8377_1_),
	   .A2 (new_n8371_),
	   .A1 (new_n8357_) );
   AOI22_X1 g1647 (
	   .ZN (new_n8377_1_),
	   .B2 (net_7220),
	   .B1 (new_n7844_),
	   .A2 (new_n8376_),
	   .A1 (new_n7837_) );
   NAND4_X1 g1646 (
	   .ZN (new_n8376_),
	   .A4 (new_n8375_),
	   .A3 (new_n8374_),
	   .A2 (new_n8373_),
	   .A1 (new_n8372_1_) );
   NAND3_X1 g1645 (
	   .ZN (new_n8375_),
	   .A3 (_net_7228),
	   .A2 (_net_7229),
	   .A1 (net_7204) );
   NAND3_X1 g1644 (
	   .ZN (new_n8374_),
	   .A3 (net_7172),
	   .A2 (_net_7229),
	   .A1 (new_n7823_) );
   NAND3_X1 g1643 (
	   .ZN (new_n8373_),
	   .A3 (_net_7228),
	   .A2 (net_7140),
	   .A1 (new_n7821_) );
   NAND2_X1 g1642 (
	   .ZN (new_n8372_1_),
	   .A2 (net_7108),
	   .A1 (new_n7819_) );
   AND3_X1 g1641 (
	   .ZN (new_n8371_),
	   .A3 (new_n8370_),
	   .A2 (new_n8369_),
	   .A1 (new_n8363_) );
   NAND2_X1 g1640 (
	   .ZN (new_n8370_),
	   .A2 (_net_6177),
	   .A1 (new_n7694_) );
   NAND2_X1 g1639 (
	   .ZN (new_n8369_),
	   .A2 (new_n7701_),
	   .A1 (new_n8368_) );
   NAND4_X1 g1638 (
	   .ZN (new_n8368_),
	   .A4 (new_n8367_1_),
	   .A3 (new_n8366_),
	   .A2 (new_n8365_),
	   .A1 (new_n8364_) );
   NAND3_X1 g1637 (
	   .ZN (new_n8367_1_),
	   .A3 (_net_7228),
	   .A2 (net_7206),
	   .A1 (_net_7229) );
   NAND3_X1 g1636 (
	   .ZN (new_n8366_),
	   .A3 (_net_7229),
	   .A2 (net_7174),
	   .A1 (new_n7823_) );
   NAND3_X1 g1635 (
	   .ZN (new_n8365_),
	   .A3 (_net_7228),
	   .A2 (net_7142),
	   .A1 (new_n7821_) );
   NAND2_X1 g1634 (
	   .ZN (new_n8364_),
	   .A2 (net_7110),
	   .A1 (new_n7819_) );
   NAND2_X1 g1633 (
	   .ZN (new_n8363_),
	   .A2 (new_n7690_),
	   .A1 (new_n8362_1_) );
   NAND4_X1 g1632 (
	   .ZN (new_n8362_1_),
	   .A4 (new_n8361_),
	   .A3 (new_n8360_),
	   .A2 (new_n8359_1_),
	   .A1 (new_n8358_) );
   NAND3_X1 g1631 (
	   .ZN (new_n8361_),
	   .A3 (_net_7228),
	   .A2 (net_7208),
	   .A1 (_net_7229) );
   NAND3_X1 g1630 (
	   .ZN (new_n8360_),
	   .A3 (net_7176),
	   .A2 (_net_7229),
	   .A1 (new_n7823_) );
   NAND3_X1 g1629 (
	   .ZN (new_n8359_1_),
	   .A3 (_net_7228),
	   .A2 (net_7144),
	   .A1 (new_n7821_) );
   NAND2_X1 g1628 (
	   .ZN (new_n8358_),
	   .A2 (net_7112),
	   .A1 (new_n7819_) );
   AND3_X1 g1627 (
	   .ZN (new_n8357_),
	   .A3 (new_n8356_),
	   .A2 (new_n8355_),
	   .A1 (new_n8354_1_) );
   NAND4_X1 g1626 (
	   .ZN (new_n8356_),
	   .A4 (new_n7678_),
	   .A3 (_net_7227),
	   .A2 (net_7188),
	   .A1 (new_n7816_) );
   NAND4_X1 g1625 (
	   .ZN (new_n8355_),
	   .A4 (new_n7683_),
	   .A3 (_net_7227),
	   .A2 (net_7124),
	   .A1 (new_n7813_) );
   NAND4_X1 g1624 (
	   .ZN (new_n8354_1_),
	   .A4 (new_n7681_1_),
	   .A3 (net_7156),
	   .A2 (_net_7227),
	   .A1 (new_n7813_) );
   CLKBUF_X1 g1623 (
	   .Z (n2189),
	   .A (_net_7813) );
   CLKBUF_X1 g1622 (
	   .Z (n2186),
	   .A (net_6443) );
   NAND4_X1 g1621 (
	   .ZN (n2177),
	   .A4 (new_n8350_1_),
	   .A3 (new_n8349_),
	   .A2 (new_n8348_),
	   .A1 (new_n8347_) );
   NAND4_X1 g1620 (
	   .ZN (new_n8350_1_),
	   .A4 (net_7708),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   NAND4_X1 g1619 (
	   .ZN (new_n8349_),
	   .A4 (new_n7364_),
	   .A3 (_net_6007),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   NAND4_X1 g1618 (
	   .ZN (new_n8348_),
	   .A4 (_net_290),
	   .A3 (x1286),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR2_X1 g1617 (
	   .ZN (new_n8347_),
	   .A2 (new_n8346_),
	   .A1 (new_n8345_1_) );
   AND2_X1 g1616 (
	   .ZN (new_n8346_),
	   .A2 (net_7737),
	   .A1 (new_n7934_) );
   NAND4_X1 g1615 (
	   .ZN (new_n8345_1_),
	   .A4 (new_n8344_),
	   .A3 (new_n8343_),
	   .A2 (new_n8342_),
	   .A1 (new_n8341_) );
   NAND4_X1 g1614 (
	   .ZN (new_n8344_),
	   .A4 (_net_173),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g1613 (
	   .ZN (new_n8343_),
	   .A3 (_net_210),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g1612 (
	   .ZN (new_n8342_),
	   .A3 (net_247),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   NAND4_X1 g1611 (
	   .ZN (new_n8341_),
	   .A4 (new_n7354_1_),
	   .A3 (net_147),
	   .A2 (x1261),
	   .A1 (new_n7370_) );
   AOI21_X1 g1610 (
	   .ZN (n2172),
	   .B2 (new_n8338_),
	   .B1 (_net_6963),
	   .A (new_n8339_) );
   OAI21_X1 g1609 (
	   .ZN (new_n8339_),
	   .B2 (_net_6963),
	   .B1 (new_n8338_),
	   .A (_net_6017) );
   AND3_X1 g1608 (
	   .ZN (new_n8338_),
	   .A3 (_net_6962),
	   .A2 (_net_5975),
	   .A1 (net_6961) );
   MUX2_X1 g1607 (
	   .Z (n2167),
	   .S (new_n7545_),
	   .B (_net_7649),
	   .A (new_n8336_) );
   OAI21_X1 g1606 (
	   .ZN (new_n8336_),
	   .B2 (new_n8335_),
	   .B1 (new_n7019_),
	   .A (new_n8334_1_) );
   INV_X1 g1605 (
	   .ZN (new_n8335_),
	   .A (net_7537) );
   AOI22_X1 g1604 (
	   .ZN (new_n8334_1_),
	   .B2 (_net_292),
	   .B1 (net_367),
	   .A2 (_net_291),
	   .A1 (net_369) );
   MUX2_X1 g1603 (
	   .Z (n2162),
	   .S (new_n7609_),
	   .B (_net_7554),
	   .A (new_n8114_) );
   CLKBUF_X1 g1602 (
	   .Z (n2157),
	   .A (_net_6140) );
   AND2_X1 g1601 (
	   .ZN (n2152),
	   .A2 (net_383),
	   .A1 (new_n7747_) );
   CLKBUF_X1 g1600 (
	   .Z (n2149),
	   .A (net_7144) );
   CLKBUF_X1 g1599 (
	   .Z (n2144),
	   .A (_net_7809) );
   OAI21_X1 g1598 (
	   .ZN (n2140),
	   .B2 (_net_7683),
	   .B1 (new_n8327_),
	   .A (new_n8324_1_) );
   NAND2_X1 g1597 (
	   .ZN (new_n8327_),
	   .A2 (new_n7262_),
	   .A1 (new_n8326_) );
   NOR2_X1 g1596 (
	   .ZN (new_n8326_),
	   .A2 (new_n8325_),
	   .A1 (new_n7024_) );
   INV_X1 g1595 (
	   .ZN (new_n8325_),
	   .A (_net_289) );
   OAI211_X1 g1594 (
	   .ZN (new_n8324_1_),
	   .C2 (new_n7024_),
	   .C1 (new_n7020_),
	   .B (_net_289),
	   .A (_net_7683) );
   CLKBUF_X1 g1593 (
	   .Z (n2136),
	   .A (net_6730) );
   CLKBUF_X1 g1592 (
	   .Z (n2132),
	   .A (net_7147) );
   CLKBUF_X1 g1591 (
	   .Z (n2127),
	   .A (_net_6114) );
   CLKBUF_X1 g1590 (
	   .Z (n2122),
	   .A (_net_7809) );
   CLKBUF_X1 g1589 (
	   .Z (n2119),
	   .A (net_6603) );
   CLKBUF_X1 g1588 (
	   .Z (n2115),
	   .A (net_6452) );
   CLKBUF_X1 g1587 (
	   .Z (n2111),
	   .A (net_7003) );
   CLKBUF_X1 g1586 (
	   .Z (n2106),
	   .A (net_6056) );
   CLKBUF_X1 g1585 (
	   .Z (n2102),
	   .A (net_6741) );
   CLKBUF_X1 g1584 (
	   .Z (n2098),
	   .A (net_6709) );
   CLKBUF_X1 g1583 (
	   .Z (n2093),
	   .A (_net_7793) );
   CLKBUF_X1 g1582 (
	   .Z (n2088),
	   .A (_net_7796) );
   NOR2_X1 g1581 (
	   .ZN (n2084),
	   .A2 (new_n8103_),
	   .A1 (new_n6952_1_) );
   CLKBUF_X1 g1580 (
	   .Z (n2079),
	   .A (_net_5968) );
   CLKBUF_X1 g1579 (
	   .Z (n2074),
	   .A (net_7799) );
   NOR3_X1 g1578 (
	   .ZN (n2070),
	   .A3 (new_n8307_1_),
	   .A2 (new_n7208_),
	   .A1 (new_n8306_) );
   AOI21_X1 g1577 (
	   .ZN (new_n8307_1_),
	   .B2 (_net_5971),
	   .B1 (net_6826),
	   .A (_net_6827) );
   NOR3_X1 g1576 (
	   .ZN (new_n8306_),
	   .A3 (new_n8305_),
	   .A2 (new_n8304_),
	   .A1 (new_n8303_1_) );
   INV_X1 g1575 (
	   .ZN (new_n8305_),
	   .A (_net_5971) );
   INV_X1 g1574 (
	   .ZN (new_n8304_),
	   .A (net_6826) );
   INV_X1 g1573 (
	   .ZN (new_n8303_1_),
	   .A (_net_6827) );
   OAI21_X1 g1572 (
	   .ZN (n2065),
	   .B2 (new_n8301_),
	   .B1 (new_n8300_),
	   .A (new_n8299_1_) );
   INV_X1 g1571 (
	   .ZN (new_n8301_),
	   .A (new_n6869_) );
   INV_X1 g1570 (
	   .ZN (new_n8300_),
	   .A (_net_6125) );
   NAND2_X1 g1569 (
	   .ZN (new_n8299_1_),
	   .A2 (new_n6854_),
	   .A1 (new_n8298_) );
   NAND2_X1 g1568 (
	   .ZN (new_n8298_),
	   .A2 (new_n8297_),
	   .A1 (new_n8296_) );
   AOI22_X1 g1567 (
	   .ZN (new_n8297_),
	   .B2 (net_6830),
	   .B1 (new_n6836_1_),
	   .A2 (net_6862),
	   .A1 (new_n6833_) );
   AOI22_X1 g1566 (
	   .ZN (new_n8296_),
	   .B2 (net_6926),
	   .B1 (new_n6873_),
	   .A2 (new_n6841_),
	   .A1 (net_6894) );
   OAI21_X1 g1565 (
	   .ZN (n2060),
	   .B2 (new_n7111_1_),
	   .B1 (new_n8294_1_),
	   .A (new_n8293_) );
   INV_X1 g1564 (
	   .ZN (new_n8294_1_),
	   .A (_net_7352) );
   NAND2_X1 g1563 (
	   .ZN (new_n8293_),
	   .A2 (new_n8292_),
	   .A1 (new_n7101_) );
   OAI221_X1 g1562 (
	   .ZN (new_n8292_),
	   .C2 (new_n7333_),
	   .C1 (new_n7106_),
	   .B2 (new_n7105_),
	   .B1 (new_n7493_),
	   .A (new_n8291_) );
   NAND2_X1 g1561 (
	   .ZN (new_n8291_),
	   .A2 (net_7240),
	   .A1 (new_n6942_) );
   OAI21_X1 g1560 (
	   .ZN (n2055),
	   .B2 (new_n6907_),
	   .B1 (new_n8289_1_),
	   .A (new_n8288_) );
   INV_X1 g1559 (
	   .ZN (new_n8289_1_),
	   .A (_net_7465) );
   NAND2_X1 g1558 (
	   .ZN (new_n8288_),
	   .A2 (new_n7874_),
	   .A1 (new_n6897_) );
   CLKBUF_X1 g1557 (
	   .Z (n2051),
	   .A (net_7391) );
   NOR2_X1 g1556 (
	   .ZN (n2046),
	   .A2 (new_n8285_),
	   .A1 (new_n8284_1_) );
   NOR3_X1 g1555 (
	   .ZN (new_n8285_),
	   .A3 (new_n7092_),
	   .A2 (new_n7077_1_),
	   .A1 (new_n7060_) );
   NOR3_X1 g1554 (
	   .ZN (new_n8284_1_),
	   .A3 (new_n7287_),
	   .A2 (_net_7093),
	   .A1 (new_n7073_) );
   OAI21_X1 g1553 (
	   .ZN (n2041),
	   .B2 (new_n6907_),
	   .B1 (new_n8282_),
	   .A (new_n8281_) );
   INV_X1 g1552 (
	   .ZN (new_n8282_),
	   .A (_net_7483) );
   NAND2_X1 g1551 (
	   .ZN (new_n8281_),
	   .A2 (new_n8280_1_),
	   .A1 (new_n6897_) );
   OAI22_X1 g1550 (
	   .ZN (new_n8280_1_),
	   .B2 (new_n6901_),
	   .B1 (new_n6903_),
	   .A2 (new_n7483_),
	   .A1 (new_n7034_) );
   CLKBUF_X1 g1549 (
	   .Z (n2036),
	   .A (net_6394) );
   CLKBUF_X1 g1548 (
	   .Z (n2031),
	   .A (_net_6122) );
   NAND2_X1 g1547 (
	   .ZN (n2026),
	   .A2 (new_n8276_1_),
	   .A1 (new_n8272_) );
   NAND2_X1 g1546 (
	   .ZN (new_n8276_1_),
	   .A2 (new_n7587_),
	   .A1 (new_n8275_) );
   NAND2_X1 g1545 (
	   .ZN (new_n8275_),
	   .A2 (new_n8274_),
	   .A1 (new_n8273_) );
   AOI22_X1 g1544 (
	   .ZN (new_n8274_),
	   .B2 (net_6695),
	   .B1 (new_n7196_),
	   .A2 (net_6727),
	   .A1 (new_n7194_1_) );
   AOI22_X1 g1543 (
	   .ZN (new_n8273_),
	   .B2 (net_6759),
	   .B1 (new_n7190_1_),
	   .A2 (new_n7188_),
	   .A1 (net_6791) );
   AOI22_X1 g1542 (
	   .ZN (new_n8272_),
	   .B2 (new_n7210_),
	   .B1 (_net_6107),
	   .A2 (new_n7203_1_),
	   .A1 (new_n8271_1_) );
   NAND2_X1 g1541 (
	   .ZN (new_n8271_1_),
	   .A2 (new_n8270_),
	   .A1 (new_n8269_) );
   AOI22_X1 g1540 (
	   .ZN (new_n8270_),
	   .B2 (net_6697),
	   .B1 (new_n7196_),
	   .A2 (net_6729),
	   .A1 (new_n7194_1_) );
   AOI22_X1 g1539 (
	   .ZN (new_n8269_),
	   .B2 (net_6761),
	   .B1 (new_n7191_),
	   .A2 (new_n7189_),
	   .A1 (net_6793) );
   OAI21_X1 g1538 (
	   .ZN (n2021),
	   .B2 (new_n8267_),
	   .B1 (new_n8266_1_),
	   .A (new_n8265_) );
   NAND2_X1 g1537 (
	   .ZN (new_n8267_),
	   .A2 (_net_6409),
	   .A1 (_net_6408) );
   OAI21_X1 g1536 (
	   .ZN (new_n8266_1_),
	   .B2 (_net_6405),
	   .B1 (_net_6406),
	   .A (_net_6407) );
   NOR2_X1 g1535 (
	   .ZN (new_n8265_),
	   .A2 (_net_6410),
	   .A1 (_net_6411) );
   AOI21_X1 g1534 (
	   .ZN (n2016),
	   .B2 (new_n7739_),
	   .B1 (new_n8263_),
	   .A (new_n8262_1_) );
   INV_X1 g1533 (
	   .ZN (new_n8263_),
	   .A (_net_7426) );
   NOR2_X1 g1532 (
	   .ZN (new_n8262_1_),
	   .A2 (n2256),
	   .A1 (new_n7739_) );
   NOR2_X1 g1531 (
	   .ZN (n2256),
	   .A2 (new_n7648_),
	   .A1 (new_n7035_) );
   CLKBUF_X1 g1530 (
	   .Z (n2011),
	   .A (_net_7818) );
   CLKBUF_X1 g1529 (
	   .Z (n2007),
	   .A (_net_7815) );
   CLKBUF_X1 g1528 (
	   .Z (n2002),
	   .A (_net_6107) );
   CLKBUF_X1 g1527 (
	   .Z (n1998),
	   .A (net_6737) );
   NOR2_X1 g1526 (
	   .ZN (n1993),
	   .A2 (new_n6933_),
	   .A1 (new_n7035_) );
   NAND4_X1 g1525 (
	   .ZN (n1988),
	   .A4 (new_n8254_),
	   .A3 (new_n8253_1_),
	   .A2 (new_n8247_),
	   .A1 (new_n8246_) );
   NAND2_X1 g1524 (
	   .ZN (new_n8254_),
	   .A2 (new_n7579_),
	   .A1 (new_n7556_) );
   AOI22_X1 g1523 (
	   .ZN (new_n8253_1_),
	   .B2 (_net_6108),
	   .B1 (new_n7210_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n8252_) );
   NAND4_X1 g1522 (
	   .ZN (new_n8252_),
	   .A4 (new_n8251_),
	   .A3 (new_n8250_),
	   .A2 (new_n8249_1_),
	   .A1 (new_n8248_) );
   NAND3_X1 g1521 (
	   .ZN (new_n8251_),
	   .A3 (_net_6824),
	   .A2 (net_6794),
	   .A1 (_net_6823) );
   NAND3_X1 g1520 (
	   .ZN (new_n8250_),
	   .A3 (_net_6824),
	   .A2 (net_6762),
	   .A1 (new_n7570_) );
   NAND3_X1 g1519 (
	   .ZN (new_n8249_1_),
	   .A3 (_net_6823),
	   .A2 (net_6730),
	   .A1 (new_n7568_) );
   NAND2_X1 g1518 (
	   .ZN (new_n8248_),
	   .A2 (net_6698),
	   .A1 (new_n7566_) );
   NAND2_X1 g1517 (
	   .ZN (new_n8247_),
	   .A2 (new_n7565_),
	   .A1 (new_n7198_) );
   NAND2_X1 g1516 (
	   .ZN (new_n8246_),
	   .A2 (new_n7587_),
	   .A1 (new_n8245_1_) );
   NAND2_X1 g1515 (
	   .ZN (new_n8245_1_),
	   .A2 (new_n8244_),
	   .A1 (new_n8243_) );
   AOI22_X1 g1514 (
	   .ZN (new_n8244_),
	   .B2 (net_6696),
	   .B1 (new_n7196_),
	   .A2 (net_6728),
	   .A1 (new_n7194_1_) );
   AOI22_X1 g1513 (
	   .ZN (new_n8243_),
	   .B2 (net_6760),
	   .B1 (new_n7191_),
	   .A2 (new_n7189_),
	   .A1 (net_6792) );
   CLKBUF_X1 g1512 (
	   .Z (n1983),
	   .A (_net_6098) );
   CLKBUF_X1 g1511 (
	   .Z (n1978),
	   .A (_net_7804) );
   CLKBUF_X1 g1510 (
	   .Z (n1973),
	   .A (_net_7803) );
   MUX2_X1 g1509 (
	   .Z (n1969),
	   .S (new_n7029_),
	   .B (_net_7594),
	   .A (new_n7806_1_) );
   CLKBUF_X1 g1508 (
	   .Z (n1964),
	   .A (_net_6150) );
   MUX2_X1 g1507 (
	   .Z (n1959),
	   .S (_net_154),
	   .B (net_325),
	   .A (_net_129) );
   CLKBUF_X1 g1506 (
	   .Z (n1954),
	   .A (_net_7817) );
   OAI21_X1 g1505 (
	   .ZN (n1950),
	   .B2 (new_n6891_),
	   .B1 (new_n8234_),
	   .A (new_n8233_) );
   INV_X1 g1504 (
	   .ZN (new_n8234_),
	   .A (new_n7951_) );
   OAI211_X1 g1503 (
	   .ZN (new_n8233_),
	   .C2 (new_n7035_),
	   .C1 (new_n7950_1_),
	   .B (_net_278),
	   .A (_net_7532) );
   OAI21_X1 g1502 (
	   .ZN (n1945),
	   .B2 (new_n6907_),
	   .B1 (new_n8231_),
	   .A (new_n8230_) );
   INV_X1 g1501 (
	   .ZN (new_n8231_),
	   .A (_net_7472) );
   NAND2_X1 g1500 (
	   .ZN (new_n8230_),
	   .A2 (new_n8229_),
	   .A1 (new_n6897_) );
   OAI221_X1 g1499 (
	   .ZN (new_n8229_),
	   .C2 (new_n6934_1_),
	   .C1 (new_n6902_1_),
	   .B2 (new_n6901_),
	   .B1 (new_n7962_1_),
	   .A (new_n8228_1_) );
   NAND2_X1 g1498 (
	   .ZN (new_n8228_1_),
	   .A2 (net_7392),
	   .A1 (new_n6898_) );
   CLKBUF_X1 g1497 (
	   .Z (n1941),
	   .A (net_6433) );
   NAND2_X1 g1496 (
	   .ZN (n1936),
	   .A2 (new_n8225_),
	   .A1 (new_n8224_1_) );
   AOI22_X1 g1495 (
	   .ZN (new_n8225_),
	   .B2 (new_n6751_),
	   .B1 (_net_7563),
	   .A2 (_net_7659),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g1494 (
	   .ZN (new_n8224_1_),
	   .B2 (_net_7627),
	   .B1 (new_n8009_),
	   .A2 (new_n6743_),
	   .A1 (_net_7595) );
   CLKBUF_X1 g1493 (
	   .Z (n1932),
	   .A (net_6995) );
   NAND2_X1 g1492 (
	   .ZN (n1927),
	   .A2 (new_n8221_),
	   .A1 (new_n8217_) );
   NAND3_X1 g1491 (
	   .ZN (new_n8221_),
	   .A3 (new_n8220_1_),
	   .A2 (new_n8219_),
	   .A1 (new_n8218_) );
   NAND2_X1 g1490 (
	   .ZN (new_n8220_1_),
	   .A2 (new_n8214_),
	   .A1 (new_n6967_) );
   INV_X1 g1489 (
	   .ZN (new_n8219_),
	   .A (new_n8215_) );
   NOR2_X1 g1488 (
	   .ZN (new_n8218_),
	   .A2 (new_n6997_),
	   .A1 (new_n6977_1_) );
   AOI22_X1 g1487 (
	   .ZN (new_n8217_),
	   .B2 (_net_6690),
	   .B1 (new_n6985_),
	   .A2 (new_n7115_),
	   .A1 (new_n8216_1_) );
   AOI22_X1 g1486 (
	   .ZN (new_n8216_1_),
	   .B2 (new_n7135_),
	   .B1 (new_n8214_),
	   .A2 (_net_6687),
	   .A1 (new_n8215_) );
   NOR2_X1 g1485 (
	   .ZN (new_n8215_),
	   .A2 (new_n8214_),
	   .A1 (new_n6967_) );
   INV_X1 g1484 (
	   .ZN (new_n8214_),
	   .A (_net_6690) );
   NAND4_X1 g1483 (
	   .ZN (n1922),
	   .A4 (new_n8212_),
	   .A3 (new_n8206_1_),
	   .A2 (new_n8204_),
	   .A1 (new_n8200_) );
   AOI22_X1 g1482 (
	   .ZN (new_n8212_),
	   .B2 (_net_6070),
	   .B1 (new_n6813_1_),
	   .A2 (new_n7166_),
	   .A1 (new_n8211_1_) );
   NAND4_X1 g1481 (
	   .ZN (new_n8211_1_),
	   .A4 (new_n8210_),
	   .A3 (new_n8209_),
	   .A2 (new_n8208_),
	   .A1 (new_n8207_) );
   NAND3_X1 g1480 (
	   .ZN (new_n8210_),
	   .A3 (_net_6554),
	   .A2 (net_6526),
	   .A1 (_net_6553) );
   NAND3_X1 g1479 (
	   .ZN (new_n8209_),
	   .A3 (net_6494),
	   .A2 (_net_6554),
	   .A1 (new_n6789_) );
   NAND3_X1 g1478 (
	   .ZN (new_n8208_),
	   .A3 (net_6462),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   NAND2_X1 g1477 (
	   .ZN (new_n8207_),
	   .A2 (net_6430),
	   .A1 (new_n6785_) );
   NAND2_X1 g1476 (
	   .ZN (new_n8206_1_),
	   .A2 (new_n6807_),
	   .A1 (new_n8205_) );
   NOR2_X1 g1475 (
	   .ZN (new_n8205_),
	   .A2 (new_n7859_),
	   .A1 (new_n6782_) );
   NAND2_X1 g1474 (
	   .ZN (new_n8204_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n8203_) );
   NAND2_X1 g1473 (
	   .ZN (new_n8203_),
	   .A2 (new_n8202_1_),
	   .A1 (new_n8201_) );
   AOI22_X1 g1472 (
	   .ZN (new_n8202_1_),
	   .B2 (net_6428),
	   .B1 (new_n6785_),
	   .A2 (net_6460),
	   .A1 (new_n6766_) );
   AOI22_X1 g1471 (
	   .ZN (new_n8201_),
	   .B2 (net_6524),
	   .B1 (new_n8139_),
	   .A2 (new_n6774_1_),
	   .A1 (net_6492) );
   NAND2_X1 g1470 (
	   .ZN (new_n8200_),
	   .A2 (new_n6784_),
	   .A1 (new_n8199_) );
   NAND2_X1 g1469 (
	   .ZN (new_n8199_),
	   .A2 (new_n8198_),
	   .A1 (new_n8197_1_) );
   AOI22_X1 g1468 (
	   .ZN (new_n8198_),
	   .B2 (net_6426),
	   .B1 (new_n6770_1_),
	   .A2 (net_6458),
	   .A1 (new_n6767_) );
   AOI22_X1 g1467 (
	   .ZN (new_n8197_1_),
	   .B2 (net_6522),
	   .B1 (new_n8139_),
	   .A2 (new_n6775_),
	   .A1 (net_6490) );
   CLKBUF_X1 g1466 (
	   .Z (n1918),
	   .A (net_7116) );
   CLKBUF_X1 g1465 (
	   .Z (n1913),
	   .A (_net_7816) );
   NOR3_X1 g1464 (
	   .ZN (n1908),
	   .A3 (new_n8193_),
	   .A2 (new_n8192_1_),
	   .A1 (new_n8191_) );
   INV_X1 g1463 (
	   .ZN (new_n8193_),
	   .A (_net_267) );
   AOI21_X1 g1462 (
	   .ZN (new_n8192_1_),
	   .B2 (_net_190),
	   .B1 (net_7378),
	   .A (_net_7379) );
   AND3_X1 g1461 (
	   .ZN (new_n8191_),
	   .A3 (_net_190),
	   .A2 (net_7378),
	   .A1 (_net_7379) );
   CLKBUF_X1 g1460 (
	   .Z (n1903),
	   .A (_net_6082) );
   NOR4_X1 g1459 (
	   .ZN (n1898),
	   .A4 (_net_6405),
	   .A3 (new_n8188_1_),
	   .A2 (new_n8187_),
	   .A1 (new_n8184_) );
   INV_X1 g1458 (
	   .ZN (new_n8188_1_),
	   .A (_net_6404) );
   NAND2_X1 g1457 (
	   .ZN (new_n8187_),
	   .A2 (new_n8186_),
	   .A1 (new_n8185_) );
   INV_X1 g1456 (
	   .ZN (new_n8186_),
	   .A (_net_6409) );
   INV_X1 g1455 (
	   .ZN (new_n8185_),
	   .A (_net_6408) );
   NAND4_X1 g1454 (
	   .ZN (new_n8184_),
	   .A4 (_net_6407),
	   .A3 (_net_6410),
	   .A2 (_net_6406),
	   .A1 (new_n8183_1_) );
   INV_X1 g1453 (
	   .ZN (new_n8183_1_),
	   .A (_net_6411) );
   NAND3_X1 g1452 (
	   .ZN (n1893),
	   .A3 (new_n8181_),
	   .A2 (new_n8174_1_),
	   .A1 (new_n8160_) );
   AOI22_X1 g1451 (
	   .ZN (new_n8181_),
	   .B2 (new_n8180_),
	   .B1 (net_7083),
	   .A2 (new_n8179_1_),
	   .A1 (new_n7060_) );
   NOR3_X2 g1450 (
	   .ZN (new_n8180_),
	   .A3 (new_n7290_),
	   .A2 (new_n8153_),
	   .A1 (new_n7067_1_) );
   NAND4_X1 g1449 (
	   .ZN (new_n8179_1_),
	   .A4 (new_n8178_),
	   .A3 (new_n8177_),
	   .A2 (new_n8176_),
	   .A1 (new_n8175_) );
   NAND3_X1 g1448 (
	   .ZN (new_n8178_),
	   .A3 (_net_7093),
	   .A2 (net_7067),
	   .A1 (_net_7094) );
   NAND3_X1 g1447 (
	   .ZN (new_n8177_),
	   .A3 (net_7035),
	   .A2 (_net_7094),
	   .A1 (new_n7048_) );
   NAND3_X1 g1446 (
	   .ZN (new_n8176_),
	   .A3 (net_7003),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   NAND2_X1 g1445 (
	   .ZN (new_n8175_),
	   .A2 (net_6971),
	   .A1 (new_n7063_) );
   AND3_X1 g1444 (
	   .ZN (new_n8174_1_),
	   .A3 (new_n8173_),
	   .A2 (new_n8172_),
	   .A1 (new_n8166_1_) );
   NAND2_X1 g1443 (
	   .ZN (new_n8173_),
	   .A2 (_net_6155),
	   .A1 (new_n7092_) );
   NAND2_X1 g1442 (
	   .ZN (new_n8172_),
	   .A2 (new_n7070_),
	   .A1 (new_n8171_) );
   NAND4_X1 g1441 (
	   .ZN (new_n8171_),
	   .A4 (new_n8170_1_),
	   .A3 (new_n8169_),
	   .A2 (new_n8168_),
	   .A1 (new_n8167_) );
   NAND3_X1 g1440 (
	   .ZN (new_n8170_1_),
	   .A3 (net_7069),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   NAND3_X1 g1439 (
	   .ZN (new_n8169_),
	   .A3 (net_7037),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g1438 (
	   .ZN (new_n8168_),
	   .A3 (net_7005),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   NAND2_X1 g1437 (
	   .ZN (new_n8167_),
	   .A2 (net_6973),
	   .A1 (new_n7063_) );
   NAND2_X1 g1436 (
	   .ZN (new_n8166_1_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n8165_) );
   NAND4_X1 g1435 (
	   .ZN (new_n8165_),
	   .A4 (new_n8164_),
	   .A3 (new_n8163_),
	   .A2 (new_n8162_),
	   .A1 (new_n8161_1_) );
   NAND3_X1 g1434 (
	   .ZN (new_n8164_),
	   .A3 (net_7071),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   NAND3_X1 g1433 (
	   .ZN (new_n8163_),
	   .A3 (net_7039),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g1432 (
	   .ZN (new_n8162_),
	   .A3 (net_7007),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   NAND2_X1 g1431 (
	   .ZN (new_n8161_1_),
	   .A2 (net_6975),
	   .A1 (new_n7063_) );
   AND3_X1 g1430 (
	   .ZN (new_n8160_),
	   .A3 (new_n8159_),
	   .A2 (new_n8157_),
	   .A1 (new_n8156_1_) );
   NAND4_X1 g1429 (
	   .ZN (new_n8159_),
	   .A4 (new_n7044_),
	   .A3 (net_7051),
	   .A2 (_net_7092),
	   .A1 (new_n8158_) );
   BUF_X4 g1428 (
	   .Z (new_n8158_),
	   .A (new_n8154_) );
   NAND4_X1 g1427 (
	   .ZN (new_n8157_),
	   .A4 (new_n7052_),
	   .A3 (net_6987),
	   .A2 (_net_7092),
	   .A1 (new_n8155_) );
   NAND4_X1 g1426 (
	   .ZN (new_n8156_1_),
	   .A4 (new_n7050_),
	   .A3 (_net_7092),
	   .A2 (net_7019),
	   .A1 (new_n8155_) );
   BUF_X4 g1425 (
	   .Z (new_n8155_),
	   .A (new_n8154_) );
   NOR2_X1 g1424 (
	   .ZN (new_n8154_),
	   .A2 (new_n8153_),
	   .A1 (new_n7067_1_) );
   INV_X1 g1423 (
	   .ZN (new_n8153_),
	   .A (new_n7057_) );
   MUX2_X1 g1422 (
	   .Z (n1888),
	   .S (new_n7504_),
	   .B (_net_7628),
	   .A (new_n8151_) );
   OAI21_X1 g1421 (
	   .ZN (new_n8151_),
	   .B2 (new_n8150_),
	   .B1 (new_n7019_),
	   .A (new_n8149_) );
   INV_X1 g1420 (
	   .ZN (new_n8150_),
	   .A (net_7548) );
   AOI22_X1 g1419 (
	   .ZN (new_n8149_),
	   .B2 (_net_291),
	   .B1 (net_380),
	   .A2 (_net_292),
	   .A1 (net_378) );
   NAND2_X1 g1418 (
	   .ZN (n1883),
	   .A2 (new_n8147_1_),
	   .A1 (new_n8143_) );
   NAND2_X1 g1417 (
	   .ZN (new_n8147_1_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n8146_) );
   NAND2_X1 g1416 (
	   .ZN (new_n8146_),
	   .A2 (new_n8145_),
	   .A1 (new_n8144_1_) );
   AOI22_X1 g1415 (
	   .ZN (new_n8145_),
	   .B2 (net_6425),
	   .B1 (new_n6770_1_),
	   .A2 (net_6457),
	   .A1 (new_n6767_) );
   AOI22_X1 g1414 (
	   .ZN (new_n8144_1_),
	   .B2 (net_6521),
	   .B1 (new_n8139_),
	   .A2 (new_n6775_),
	   .A1 (net_6489) );
   AOI22_X1 g1413 (
	   .ZN (new_n8143_),
	   .B2 (new_n6813_1_),
	   .B1 (_net_6067),
	   .A2 (new_n7166_),
	   .A1 (new_n8142_) );
   NAND2_X1 g1412 (
	   .ZN (new_n8142_),
	   .A2 (new_n8141_),
	   .A1 (new_n8140_1_) );
   AOI22_X1 g1411 (
	   .ZN (new_n8141_),
	   .B2 (net_6427),
	   .B1 (new_n6770_1_),
	   .A2 (net_6459),
	   .A1 (new_n6767_) );
   AOI22_X1 g1410 (
	   .ZN (new_n8140_1_),
	   .B2 (net_6523),
	   .B1 (new_n8139_),
	   .A2 (new_n6775_),
	   .A1 (net_6491) );
   INV_X1 g1409 (
	   .ZN (new_n8139_),
	   .A (new_n7856_) );
   MUX2_X1 g1408 (
	   .Z (n1878),
	   .S (new_n7029_),
	   .B (_net_7600),
	   .A (new_n7501_1_) );
   CLKBUF_X1 g1407 (
	   .Z (n1874),
	   .A (net_6599) );
   OAI21_X1 g1406 (
	   .ZN (n1869),
	   .B2 (new_n6957_1_),
	   .B1 (new_n8135_1_),
	   .A (new_n8134_) );
   INV_X1 g1405 (
	   .ZN (new_n8135_1_),
	   .A (_net_7255) );
   NAND2_X1 g1404 (
	   .ZN (new_n8134_),
	   .A2 (new_n8133_),
	   .A1 (new_n6949_) );
   OAI221_X1 g1403 (
	   .ZN (new_n8133_),
	   .C2 (new_n8132_),
	   .C1 (new_n7105_),
	   .B2 (new_n7106_),
	   .B1 (new_n7666_1_),
	   .A (new_n8131_) );
   INV_X1 g1402 (
	   .ZN (new_n8132_),
	   .A (net_333) );
   NAND2_X1 g1401 (
	   .ZN (new_n8131_),
	   .A2 (net_7239),
	   .A1 (new_n6942_) );
   CLKBUF_X1 g1400 (
	   .Z (n1865),
	   .A (net_6699) );
   AND2_X1 g1399 (
	   .ZN (n1860),
	   .A2 (net_153),
	   .A1 (_net_7768) );
   CLKBUF_X1 g1398 (
	   .Z (n1855),
	   .A (x1382) );
   AND2_X1 g1397 (
	   .ZN (n1851),
	   .A2 (_net_6222),
	   .A1 (new_n7239_) );
   AND2_X1 g1396 (
	   .ZN (n1846),
	   .A2 (_net_6291),
	   .A1 (new_n7239_) );
   NAND2_X1 g1395 (
	   .ZN (n1841),
	   .A2 (new_n8124_),
	   .A1 (new_n8120_) );
   NAND2_X1 g1394 (
	   .ZN (new_n8124_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n8123_) );
   NAND2_X1 g1393 (
	   .ZN (new_n8123_),
	   .A2 (new_n8122_),
	   .A1 (new_n8121_1_) );
   AOI22_X1 g1392 (
	   .ZN (new_n8122_),
	   .B2 (net_6560),
	   .B1 (new_n6990_1_),
	   .A2 (net_6592),
	   .A1 (new_n6971_) );
   AOI22_X1 g1391 (
	   .ZN (new_n8121_1_),
	   .B2 (net_6656),
	   .B1 (new_n6968_),
	   .A2 (new_n6966_),
	   .A1 (net_6624) );
   AOI22_X1 g1390 (
	   .ZN (new_n8120_),
	   .B2 (new_n6985_),
	   .B1 (_net_6087),
	   .A2 (new_n6980_),
	   .A1 (new_n8119_) );
   NAND2_X1 g1389 (
	   .ZN (new_n8119_),
	   .A2 (new_n8118_),
	   .A1 (new_n8117_) );
   AOI22_X1 g1388 (
	   .ZN (new_n8118_),
	   .B2 (net_6562),
	   .B1 (new_n6990_1_),
	   .A2 (net_6594),
	   .A1 (new_n6989_) );
   AOI22_X1 g1387 (
	   .ZN (new_n8117_),
	   .B2 (net_6658),
	   .B1 (new_n6968_),
	   .A2 (new_n6987_),
	   .A1 (net_6626) );
   CLKBUF_X1 g1386 (
	   .Z (n1836),
	   .A (x1432) );
   MUX2_X1 g1385 (
	   .Z (n1832),
	   .S (new_n7545_),
	   .B (_net_7650),
	   .A (new_n8114_) );
   OAI21_X1 g1384 (
	   .ZN (new_n8114_),
	   .B2 (new_n8113_),
	   .B1 (new_n7020_),
	   .A (new_n8112_1_) );
   INV_X1 g1383 (
	   .ZN (new_n8113_),
	   .A (net_7538) );
   AOI22_X1 g1382 (
	   .ZN (new_n8112_1_),
	   .B2 (net_368),
	   .B1 (_net_292),
	   .A2 (net_370),
	   .A1 (_net_291) );
   CLKBUF_X1 g1381 (
	   .Z (n1827),
	   .A (_net_6072) );
   CLKBUF_X1 g1380 (
	   .Z (n1822),
	   .A (_net_6093) );
   CLKBUF_X1 g1379 (
	   .Z (n1817),
	   .A (_net_6175) );
   OAI21_X1 g1378 (
	   .ZN (n1812),
	   .B2 (new_n7111_1_),
	   .B1 (new_n8107_1_),
	   .A (new_n8106_) );
   INV_X1 g1377 (
	   .ZN (new_n8107_1_),
	   .A (_net_7359) );
   NAND2_X1 g1376 (
	   .ZN (new_n8106_),
	   .A2 (new_n8105_),
	   .A1 (new_n7101_) );
   OAI221_X1 g1375 (
	   .ZN (new_n8105_),
	   .C2 (new_n8104_),
	   .C1 (new_n7105_),
	   .B2 (new_n7106_),
	   .B1 (new_n8103_),
	   .A (new_n8102_1_) );
   INV_X1 g1374 (
	   .ZN (new_n8104_),
	   .A (net_341) );
   INV_X1 g1373 (
	   .ZN (new_n8103_),
	   .A (net_339) );
   NAND2_X1 g1372 (
	   .ZN (new_n8102_1_),
	   .A2 (net_7247),
	   .A1 (new_n6942_) );
   OAI21_X1 g1371 (
	   .ZN (n1807),
	   .B2 (new_n7225_),
	   .B1 (new_n8100_),
	   .A (new_n8099_) );
   INV_X1 g1370 (
	   .ZN (new_n8100_),
	   .A (_net_7328) );
   NAND2_X1 g1369 (
	   .ZN (new_n8099_),
	   .A2 (new_n7531_),
	   .A1 (new_n7222_) );
   AND2_X1 g1368 (
	   .ZN (n1802),
	   .A2 (_net_6219),
	   .A1 (new_n7239_) );
   CLKBUF_X1 g1367 (
	   .Z (n1797),
	   .A (_net_6120) );
   AND2_X1 g1366 (
	   .ZN (n1787),
	   .A2 (_net_6295),
	   .A1 (new_n7239_) );
   CLKBUF_X1 g1365 (
	   .Z (n1782),
	   .A (_net_7800) );
   CLKBUF_X1 g1364 (
	   .Z (n1779),
	   .A (net_7551) );
   CLKBUF_X1 g1363 (
	   .Z (n1775),
	   .A (net_6602) );
   OAI21_X1 g1362 (
	   .ZN (n1770),
	   .B2 (new_n7437_1_),
	   .B1 (new_n8091_),
	   .A (new_n8090_) );
   INV_X1 g1361 (
	   .ZN (new_n8091_),
	   .A (_net_7794) );
   NAND2_X1 g1360 (
	   .ZN (new_n8090_),
	   .A2 (_net_5985),
	   .A1 (new_n7437_1_) );
   CLKBUF_X1 g1359 (
	   .Z (n1765),
	   .A (_net_7821) );
   CLKBUF_X1 g1358 (
	   .Z (n1761),
	   .A (net_6570) );
   CLKBUF_X1 g1357 (
	   .Z (n1756),
	   .A (_net_7796) );
   NOR2_X1 g1356 (
	   .ZN (n1752),
	   .A2 (new_n6903_),
	   .A1 (new_n7035_) );
   NAND3_X1 g1355 (
	   .ZN (n1747),
	   .A3 (new_n8084_),
	   .A2 (new_n8080_1_),
	   .A1 (new_n8074_) );
   AND3_X1 g1354 (
	   .ZN (new_n8084_),
	   .A3 (new_n8083_),
	   .A2 (new_n8082_),
	   .A1 (new_n8081_) );
   NAND2_X1 g1353 (
	   .ZN (new_n8083_),
	   .A2 (_net_6077),
	   .A1 (new_n6813_1_) );
   NAND2_X1 g1352 (
	   .ZN (new_n8082_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n7159_) );
   NAND2_X1 g1351 (
	   .ZN (new_n8081_),
	   .A2 (new_n7166_),
	   .A1 (new_n7172_1_) );
   AOI22_X1 g1350 (
	   .ZN (new_n8080_1_),
	   .B2 (new_n8079_),
	   .B1 (new_n6784_),
	   .A2 (new_n6779_1_),
	   .A1 (net_6545) );
   NAND4_X1 g1349 (
	   .ZN (new_n8079_),
	   .A4 (new_n8078_),
	   .A3 (new_n8077_),
	   .A2 (new_n8076_),
	   .A1 (new_n8075_1_) );
   NAND3_X1 g1348 (
	   .ZN (new_n8078_),
	   .A3 (net_6529),
	   .A2 (_net_6554),
	   .A1 (_net_6553) );
   NAND3_X1 g1347 (
	   .ZN (new_n8077_),
	   .A3 (_net_6554),
	   .A2 (net_6497),
	   .A1 (new_n6789_) );
   NAND3_X1 g1346 (
	   .ZN (new_n8076_),
	   .A3 (net_6465),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   NAND2_X1 g1345 (
	   .ZN (new_n8075_1_),
	   .A2 (net_6433),
	   .A1 (new_n6785_) );
   AND3_X1 g1344 (
	   .ZN (new_n8074_),
	   .A3 (new_n8073_),
	   .A2 (new_n8072_1_),
	   .A1 (new_n8071_) );
   NAND4_X1 g1343 (
	   .ZN (new_n8073_),
	   .A4 (new_n6775_),
	   .A3 (_net_6552),
	   .A2 (net_6513),
	   .A1 (new_n6772_) );
   NAND4_X1 g1342 (
	   .ZN (new_n8072_1_),
	   .A4 (new_n6770_1_),
	   .A3 (_net_6552),
	   .A2 (net_6449),
	   .A1 (new_n6764_) );
   NAND4_X1 g1341 (
	   .ZN (new_n8071_),
	   .A4 (new_n6767_),
	   .A3 (_net_6552),
	   .A2 (net_6481),
	   .A1 (new_n6764_) );
   MUX2_X1 g1340 (
	   .Z (n1742),
	   .S (new_n7437_1_),
	   .B (_net_5996),
	   .A (net_7802) );
   OAI21_X1 g1339 (
	   .ZN (n1737),
	   .B2 (new_n6907_),
	   .B1 (new_n8068_),
	   .A (new_n8067_1_) );
   INV_X1 g1338 (
	   .ZN (new_n8068_),
	   .A (_net_7468) );
   NAND2_X1 g1337 (
	   .ZN (new_n8067_1_),
	   .A2 (new_n8066_),
	   .A1 (new_n6897_) );
   OAI21_X1 g1336 (
	   .ZN (new_n8066_),
	   .B2 (new_n8065_),
	   .B1 (new_n7034_),
	   .A (new_n8064_1_) );
   INV_X1 g1335 (
	   .ZN (new_n8065_),
	   .A (net_7388) );
   AOI22_X1 g1334 (
	   .ZN (new_n8064_1_),
	   .B2 (_net_281),
	   .B1 (net_349),
	   .A2 (_net_280),
	   .A1 (net_351) );
   CLKBUF_X1 g1333 (
	   .Z (n1732),
	   .A (_net_7809) );
   NAND3_X1 g1332 (
	   .ZN (n1727),
	   .A3 (new_n8061_),
	   .A2 (new_n8055_),
	   .A1 (new_n8051_1_) );
   AOI22_X1 g1331 (
	   .ZN (new_n8061_),
	   .B2 (net_7223),
	   .B1 (new_n7844_),
	   .A2 (new_n8060_),
	   .A1 (new_n7837_) );
   NAND4_X1 g1330 (
	   .ZN (new_n8060_),
	   .A4 (new_n8059_1_),
	   .A3 (new_n8058_),
	   .A2 (new_n8057_),
	   .A1 (new_n8056_1_) );
   NAND3_X1 g1329 (
	   .ZN (new_n8059_1_),
	   .A3 (_net_7228),
	   .A2 (net_7207),
	   .A1 (_net_7229) );
   NAND3_X1 g1328 (
	   .ZN (new_n8058_),
	   .A3 (net_7175),
	   .A2 (_net_7229),
	   .A1 (new_n7823_) );
   NAND3_X1 g1327 (
	   .ZN (new_n8057_),
	   .A3 (net_7143),
	   .A2 (_net_7228),
	   .A1 (new_n7821_) );
   NAND2_X1 g1326 (
	   .ZN (new_n8056_1_),
	   .A2 (net_7111),
	   .A1 (new_n7819_) );
   AND3_X1 g1325 (
	   .ZN (new_n8055_),
	   .A3 (new_n8054_),
	   .A2 (new_n8053_),
	   .A1 (new_n8052_) );
   NAND2_X1 g1324 (
	   .ZN (new_n8054_),
	   .A2 (_net_6180),
	   .A1 (new_n7694_) );
   NAND2_X1 g1323 (
	   .ZN (new_n8053_),
	   .A2 (new_n7701_),
	   .A1 (new_n7842_) );
   NAND2_X1 g1322 (
	   .ZN (new_n8052_),
	   .A2 (new_n7690_),
	   .A1 (new_n7826_1_) );
   AND3_X1 g1321 (
	   .ZN (new_n8051_1_),
	   .A3 (new_n8050_),
	   .A2 (new_n8049_),
	   .A1 (new_n8048_) );
   NAND4_X1 g1320 (
	   .ZN (new_n8050_),
	   .A4 (new_n7678_),
	   .A3 (_net_7227),
	   .A2 (net_7191),
	   .A1 (new_n7816_) );
   NAND4_X1 g1319 (
	   .ZN (new_n8049_),
	   .A4 (new_n7683_),
	   .A3 (net_7127),
	   .A2 (_net_7227),
	   .A1 (new_n7813_) );
   NAND4_X1 g1318 (
	   .ZN (new_n8048_),
	   .A4 (new_n7681_1_),
	   .A3 (_net_7227),
	   .A2 (net_7159),
	   .A1 (new_n7813_) );
   CLKBUF_X1 g1317 (
	   .Z (n1722),
	   .A (_net_7818) );
   CLKBUF_X1 g1316 (
	   .Z (n1718),
	   .A (_net_7803) );
   OAI21_X1 g1315 (
	   .ZN (n1714),
	   .B2 (new_n7111_1_),
	   .B1 (new_n8044_),
	   .A (new_n8043_) );
   INV_X1 g1314 (
	   .ZN (new_n8044_),
	   .A (_net_7358) );
   NAND2_X1 g1313 (
	   .ZN (new_n8043_),
	   .A2 (new_n8042_1_),
	   .A1 (new_n7101_) );
   OAI21_X1 g1312 (
	   .ZN (new_n8042_1_),
	   .B2 (new_n8041_),
	   .B1 (new_n6951_),
	   .A (new_n8040_) );
   INV_X1 g1311 (
	   .ZN (new_n8041_),
	   .A (net_7246) );
   AOI22_X1 g1310 (
	   .ZN (new_n8040_),
	   .B2 (net_340),
	   .B1 (_net_269),
	   .A2 (net_338),
	   .A1 (_net_270) );
   CLKBUF_X1 g1309 (
	   .Z (n1709),
	   .A (_net_7800) );
   CLKBUF_X1 g1308 (
	   .Z (n1704),
	   .A (_net_7805) );
   CLKBUF_X1 g1307 (
	   .Z (n1701),
	   .A (net_6432) );
   NAND4_X1 g1306 (
	   .ZN (n1696),
	   .A4 (new_n8035_),
	   .A3 (new_n8031_),
	   .A2 (new_n8027_),
	   .A1 (new_n8023_) );
   NAND2_X1 g1305 (
	   .ZN (new_n8035_),
	   .A2 (new_n7837_),
	   .A1 (new_n8034_) );
   NAND2_X1 g1304 (
	   .ZN (new_n8034_),
	   .A2 (new_n8033_1_),
	   .A1 (new_n8032_) );
   AOI22_X1 g1303 (
	   .ZN (new_n8033_1_),
	   .B2 (net_7099),
	   .B1 (new_n7683_),
	   .A2 (net_7131),
	   .A1 (new_n7680_) );
   AOI22_X1 g1302 (
	   .ZN (new_n8032_),
	   .B2 (net_7163),
	   .B1 (new_n7677_),
	   .A2 (new_n7676_1_),
	   .A1 (net_7195) );
   NAND2_X1 g1301 (
	   .ZN (new_n8031_),
	   .A2 (new_n7701_),
	   .A1 (new_n8030_) );
   NAND2_X1 g1300 (
	   .ZN (new_n8030_),
	   .A2 (new_n8029_),
	   .A1 (new_n8028_1_) );
   AOI22_X1 g1299 (
	   .ZN (new_n8029_),
	   .B2 (net_7101),
	   .B1 (new_n7683_),
	   .A2 (net_7133),
	   .A1 (new_n7681_1_) );
   AOI22_X1 g1298 (
	   .ZN (new_n8028_1_),
	   .B2 (net_7165),
	   .B1 (new_n7678_),
	   .A2 (new_n7676_1_),
	   .A1 (net_7197) );
   NAND2_X1 g1297 (
	   .ZN (new_n8027_),
	   .A2 (new_n7826_1_),
	   .A1 (new_n8026_) );
   NOR2_X1 g1296 (
	   .ZN (new_n8026_),
	   .A2 (new_n8025_),
	   .A1 (new_n8024_1_) );
   INV_X1 g1295 (
	   .ZN (new_n8025_),
	   .A (_net_7227) );
   INV_X1 g1294 (
	   .ZN (new_n8024_1_),
	   .A (new_n7812_) );
   AOI22_X1 g1293 (
	   .ZN (new_n8023_),
	   .B2 (new_n7694_),
	   .B1 (_net_6168),
	   .A2 (new_n7690_),
	   .A1 (new_n8022_) );
   NAND2_X1 g1292 (
	   .ZN (new_n8022_),
	   .A2 (new_n8021_),
	   .A1 (new_n8020_) );
   AOI22_X1 g1291 (
	   .ZN (new_n8021_),
	   .B2 (net_7103),
	   .B1 (new_n7819_),
	   .A2 (net_7135),
	   .A1 (new_n7680_) );
   AOI22_X1 g1290 (
	   .ZN (new_n8020_),
	   .B2 (net_7167),
	   .B1 (new_n7677_),
	   .A2 (new_n7676_1_),
	   .A1 (net_7199) );
   CLKBUF_X1 g1289 (
	   .Z (n1691),
	   .A (_net_7805) );
   CLKBUF_X1 g1288 (
	   .Z (n1686),
	   .A (_net_7817) );
   CLKBUF_X1 g1287 (
	   .Z (n1681),
	   .A (_net_7824) );
   MUX2_X1 g1286 (
	   .Z (n1677),
	   .S (new_n6823_),
	   .B (_net_6042),
	   .A (_net_7804) );
   CLKBUF_X1 g1285 (
	   .Z (n1673),
	   .A (net_6723) );
   CLKBUF_X1 g1284 (
	   .Z (n1668),
	   .A (_net_5980) );
   CLKBUF_X1 g1283 (
	   .Z (n1663),
	   .A (net_6061) );
   NAND2_X1 g1282 (
	   .ZN (n1658),
	   .A2 (new_n8011_),
	   .A1 (new_n8010_1_) );
   AOI22_X1 g1281 (
	   .ZN (new_n8011_),
	   .B2 (new_n6751_),
	   .B1 (_net_7567),
	   .A2 (_net_7663),
	   .A1 (new_n6749_1_) );
   AOI22_X1 g1280 (
	   .ZN (new_n8010_1_),
	   .B2 (_net_7631),
	   .B1 (new_n8009_),
	   .A2 (new_n6743_),
	   .A1 (_net_7599) );
   BUF_X4 g1279 (
	   .Z (new_n8009_),
	   .A (new_n6745_) );
   CLKBUF_X1 g1278 (
	   .Z (n1653),
	   .A (net_135) );
   CLKBUF_X1 g1277 (
	   .Z (n1649),
	   .A (net_7124) );
   NAND2_X1 g1276 (
	   .ZN (n1644),
	   .A2 (new_n8005_1_),
	   .A1 (new_n8004_) );
   AOI22_X1 g1275 (
	   .ZN (new_n8005_1_),
	   .B2 (_net_7582),
	   .B1 (new_n6755_),
	   .A2 (net_7614),
	   .A1 (new_n6743_) );
   AOI22_X1 g1274 (
	   .ZN (new_n8004_),
	   .B2 (net_7646),
	   .B1 (new_n6746_1_),
	   .A2 (new_n7970_1_),
	   .A1 (net_7678) );
   AND2_X1 g1273 (
	   .ZN (n1639),
	   .A2 (net_340),
	   .A1 (new_n7102_1_) );
   MUX2_X1 g1272 (
	   .Z (n1634),
	   .S (new_n7609_),
	   .B (_net_7570),
	   .A (new_n8001_) );
   OAI21_X1 g1271 (
	   .ZN (new_n8001_),
	   .B2 (new_n8000_),
	   .B1 (new_n7215_),
	   .A (new_n7999_) );
   INV_X1 g1270 (
	   .ZN (new_n8000_),
	   .A (net_384) );
   NAND2_X1 g1269 (
	   .ZN (new_n7999_),
	   .A2 (net_372),
	   .A1 (new_n7018_1_) );
   CLKBUF_X1 g1268 (
	   .Z (n1629),
	   .A (_net_7810) );
   MUX2_X1 g1267 (
	   .Z (n1624),
	   .S (new_n7285_),
	   .B (_net_7696),
	   .A (_net_7798) );
   CLKBUF_X1 g1266 (
	   .Z (n1619),
	   .A (_net_7796) );
   CLKBUF_X1 g1265 (
	   .Z (n1615),
	   .A (_net_7814) );
   OAI21_X1 g1264 (
	   .ZN (n1610),
	   .B2 (new_n7736_),
	   .B1 (new_n7993_),
	   .A (new_n7992_) );
   INV_X1 g1263 (
	   .ZN (new_n7993_),
	   .A (_net_7498) );
   NAND2_X1 g1262 (
	   .ZN (new_n7992_),
	   .A2 (new_n7991_),
	   .A1 (new_n7733_) );
   OAI21_X1 g1261 (
	   .ZN (new_n7991_),
	   .B2 (new_n7990_),
	   .B1 (new_n7034_),
	   .A (new_n7989_1_) );
   INV_X1 g1260 (
	   .ZN (new_n7990_),
	   .A (net_7386) );
   AOI22_X1 g1259 (
	   .ZN (new_n7989_1_),
	   .B2 (net_349),
	   .B1 (_net_280),
	   .A2 (_net_281),
	   .A1 (net_347) );
   OAI221_X1 g1258 (
	   .ZN (n1605),
	   .C2 (new_n7312_1_),
	   .C1 (new_n7987_),
	   .B2 (new_n7986_),
	   .B1 (new_n7110_),
	   .A (new_n7985_1_) );
   INV_X1 g1257 (
	   .ZN (new_n7987_),
	   .A (_net_7291) );
   BUF_X4 g1256 (
	   .Z (new_n7986_),
	   .A (new_n6919_1_) );
   AOI22_X1 g1255 (
	   .ZN (new_n7985_1_),
	   .B2 (_net_7259),
	   .B1 (new_n6913_),
	   .A2 (_net_7323),
	   .A1 (new_n6911_) );
   INV_X1 g1254 (
	   .ZN (n1600),
	   .A (new_n7983_) );
   NAND2_X1 g1253 (
	   .ZN (new_n7983_),
	   .A2 (net_6056),
	   .A1 (_net_7791) );
   CLKBUF_X1 g1252 (
	   .Z (n1596),
	   .A (net_6732) );
   CLKBUF_X1 g1251 (
	   .Z (n1591),
	   .A (net_6387) );
   CLKBUF_X1 g1250 (
	   .Z (n1587),
	   .A (net_6584) );
   OAI221_X1 g1249 (
	   .ZN (n1582),
	   .C2 (new_n7978_),
	   .C1 (new_n7956_),
	   .B2 (new_n7955_1_),
	   .B1 (new_n7977_),
	   .A (new_n7976_) );
   XNOR2_X1 g1248 (
	   .ZN (new_n7978_),
	   .B (_net_7535),
	   .A (new_n7730_) );
   INV_X1 g1247 (
	   .ZN (new_n7977_),
	   .A (_net_7535) );
   NAND3_X1 g1246 (
	   .ZN (new_n7976_),
	   .A3 (new_n7975_1_),
	   .A2 (new_n6898_),
	   .A1 (new_n7951_) );
   XNOR2_X1 g1245 (
	   .ZN (new_n7975_1_),
	   .B (_net_7535),
	   .A (new_n7953_) );
   CLKBUF_X1 g1244 (
	   .Z (n1577),
	   .A (net_6388) );
   NAND2_X1 g1243 (
	   .ZN (n1572),
	   .A2 (new_n7972_),
	   .A1 (new_n7971_) );
   AOI22_X1 g1242 (
	   .ZN (new_n7972_),
	   .B2 (_net_7580),
	   .B1 (new_n6755_),
	   .A2 (net_7612),
	   .A1 (new_n6743_) );
   AOI22_X1 g1241 (
	   .ZN (new_n7971_),
	   .B2 (net_7644),
	   .B1 (new_n6746_1_),
	   .A2 (new_n7970_1_),
	   .A1 (net_7676) );
   BUF_X4 g1240 (
	   .Z (new_n7970_1_),
	   .A (new_n6748_) );
   CLKBUF_X1 g1239 (
	   .Z (n1568),
	   .A (net_6888) );
   CLKBUF_X1 g1238 (
	   .Z (n1564),
	   .A (net_6482) );
   CLKBUF_X1 g1237 (
	   .Z (n1560),
	   .A (net_7126) );
   OAI21_X1 g1236 (
	   .ZN (n1555),
	   .B2 (new_n7652_),
	   .B1 (new_n7965_),
	   .A (new_n7964_) );
   INV_X1 g1235 (
	   .ZN (new_n7965_),
	   .A (_net_7406) );
   NAND2_X1 g1234 (
	   .ZN (new_n7964_),
	   .A2 (new_n7963_),
	   .A1 (new_n7646_) );
   OAI221_X1 g1233 (
	   .ZN (new_n7963_),
	   .C2 (new_n6902_1_),
	   .C1 (new_n7962_1_),
	   .B2 (new_n6901_),
	   .B1 (new_n7961_),
	   .A (new_n7960_) );
   INV_X1 g1232 (
	   .ZN (new_n7962_1_),
	   .A (net_353) );
   INV_X1 g1231 (
	   .ZN (new_n7961_),
	   .A (net_351) );
   NAND2_X1 g1230 (
	   .ZN (new_n7960_),
	   .A2 (net_7390),
	   .A1 (new_n6898_) );
   CLKBUF_X1 g1229 (
	   .Z (n1551),
	   .A (net_7146) );
   OAI221_X1 g1228 (
	   .ZN (n1546),
	   .C2 (new_n7957_),
	   .C1 (new_n7956_),
	   .B2 (new_n7955_1_),
	   .B1 (new_n6893_),
	   .A (new_n7954_) );
   NOR2_X1 g1227 (
	   .ZN (new_n7957_),
	   .A2 (new_n7269_),
	   .A1 (new_n6894_) );
   NAND2_X1 g1226 (
	   .ZN (new_n7956_),
	   .A2 (new_n7035_),
	   .A1 (new_n7951_) );
   NAND2_X1 g1225 (
	   .ZN (new_n7955_1_),
	   .A2 (_net_278),
	   .A1 (new_n7950_1_) );
   NAND4_X1 g1224 (
	   .ZN (new_n7954_),
	   .A4 (new_n7953_),
	   .A3 (new_n7952_),
	   .A2 (new_n6898_),
	   .A1 (new_n7951_) );
   NAND3_X1 g1223 (
	   .ZN (new_n7953_),
	   .A3 (_net_7533),
	   .A2 (_net_7532),
	   .A1 (_net_7534) );
   OAI21_X1 g1222 (
	   .ZN (new_n7952_),
	   .B2 (new_n7268_),
	   .B1 (new_n6890_1_),
	   .A (new_n6893_) );
   NOR2_X1 g1221 (
	   .ZN (new_n7951_),
	   .A2 (new_n7508_),
	   .A1 (new_n7950_1_) );
   NAND2_X1 g1220 (
	   .ZN (new_n7950_1_),
	   .A2 (new_n7949_),
	   .A1 (n2181) );
   INV_X1 g1219 (
	   .ZN (new_n7949_),
	   .A (_net_7763) );
   NOR2_X1 g1218 (
	   .ZN (n2181),
	   .A2 (new_n6887_),
	   .A1 (new_n6886_1_) );
   NAND4_X1 g1217 (
	   .ZN (n1542),
	   .A4 (new_n7946_),
	   .A3 (new_n7944_),
	   .A2 (new_n7943_),
	   .A1 (new_n7942_1_) );
   NAND4_X1 g1216 (
	   .ZN (new_n7946_),
	   .A4 (new_n7364_),
	   .A3 (net_6013),
	   .A2 (x1322),
	   .A1 (new_n7945_1_) );
   BUF_X4 g1215 (
	   .Z (new_n7945_1_),
	   .A (new_n7399_) );
   NAND4_X1 g1214 (
	   .ZN (new_n7944_),
	   .A4 (net_296),
	   .A3 (x1286),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NAND4_X1 g1213 (
	   .ZN (new_n7943_),
	   .A4 (net_7714),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR3_X1 g1212 (
	   .ZN (new_n7942_1_),
	   .A3 (new_n7941_),
	   .A2 (new_n7940_),
	   .A1 (new_n7935_) );
   AND3_X1 g1211 (
	   .ZN (new_n7941_),
	   .A3 (new_n7382_),
	   .A2 (net_253),
	   .A1 (new_n7381_1_) );
   OAI22_X1 g1210 (
	   .ZN (new_n7940_),
	   .B2 (new_n7939_),
	   .B1 (new_n7938_),
	   .A2 (new_n7937_1_),
	   .A1 (new_n7936_) );
   INV_X1 g1209 (
	   .ZN (new_n7939_),
	   .A (net_179) );
   NAND3_X1 g1208 (
	   .ZN (new_n7938_),
	   .A3 (x1231),
	   .A2 (new_n7394_),
	   .A1 (new_n7392_) );
   INV_X1 g1207 (
	   .ZN (new_n7937_1_),
	   .A (net_216) );
   NAND2_X2 g1206 (
	   .ZN (new_n7936_),
	   .A2 (new_n7388_),
	   .A1 (new_n7386_1_) );
   AND2_X1 g1205 (
	   .ZN (new_n7935_),
	   .A2 (net_7743),
	   .A1 (new_n7934_) );
   INV_X1 g1204 (
	   .ZN (new_n7934_),
	   .A (new_n7377_) );
   CLKBUF_X1 g1203 (
	   .Z (n1538),
	   .A (net_7247) );
   OAI221_X1 g1202 (
	   .ZN (n1533),
	   .C2 (new_n7306_),
	   .C1 (new_n7931_),
	   .B2 (new_n7303_),
	   .B1 (new_n7930_),
	   .A (new_n7929_1_) );
   INV_X1 g1201 (
	   .ZN (new_n7931_),
	   .A (_net_7507) );
   INV_X1 g1200 (
	   .ZN (new_n7930_),
	   .A (_net_7475) );
   AOI22_X1 g1199 (
	   .ZN (new_n7929_1_),
	   .B2 (_net_7411),
	   .B1 (new_n7298_),
	   .A2 (_net_7443),
	   .A1 (new_n7296_) );
   CLKBUF_X1 g1198 (
	   .Z (n1528),
	   .A (_net_6179) );
   CLKBUF_X1 g1197 (
	   .Z (n1524),
	   .A (net_7106) );
   NAND3_X1 g1196 (
	   .ZN (n1519),
	   .A3 (new_n7925_),
	   .A2 (new_n7919_),
	   .A1 (new_n7905_) );
   AOI22_X1 g1195 (
	   .ZN (new_n7925_),
	   .B2 (new_n7136_),
	   .B1 (net_6678),
	   .A2 (new_n7924_1_),
	   .A1 (new_n7013_1_) );
   NAND4_X1 g1194 (
	   .ZN (new_n7924_1_),
	   .A4 (new_n7923_),
	   .A3 (new_n7922_),
	   .A2 (new_n7921_),
	   .A1 (new_n7920_1_) );
   NAND3_X1 g1193 (
	   .ZN (new_n7923_),
	   .A3 (net_6662),
	   .A2 (_net_6689),
	   .A1 (_net_6688) );
   NAND3_X1 g1192 (
	   .ZN (new_n7922_),
	   .A3 (net_6630),
	   .A2 (_net_6689),
	   .A1 (new_n7004_) );
   NAND3_X1 g1191 (
	   .ZN (new_n7921_),
	   .A3 (net_6598),
	   .A2 (_net_6688),
	   .A1 (new_n7002_) );
   NAND2_X1 g1190 (
	   .ZN (new_n7920_1_),
	   .A2 (net_6566),
	   .A1 (new_n6973_) );
   AND3_X1 g1189 (
	   .ZN (new_n7919_),
	   .A3 (new_n7918_),
	   .A2 (new_n7917_),
	   .A1 (new_n7911_1_) );
   NAND2_X1 g1188 (
	   .ZN (new_n7918_),
	   .A2 (_net_6095),
	   .A1 (new_n6985_) );
   NAND2_X1 g1187 (
	   .ZN (new_n7917_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n7916_1_) );
   NAND4_X1 g1186 (
	   .ZN (new_n7916_1_),
	   .A4 (new_n7915_),
	   .A3 (new_n7914_),
	   .A2 (new_n7913_),
	   .A1 (new_n7912_) );
   NAND3_X1 g1185 (
	   .ZN (new_n7915_),
	   .A3 (_net_6689),
	   .A2 (_net_6688),
	   .A1 (net_6664) );
   NAND3_X1 g1184 (
	   .ZN (new_n7914_),
	   .A3 (_net_6689),
	   .A2 (net_6632),
	   .A1 (new_n7004_) );
   NAND3_X1 g1183 (
	   .ZN (new_n7913_),
	   .A3 (net_6600),
	   .A2 (_net_6688),
	   .A1 (new_n7002_) );
   NAND2_X1 g1182 (
	   .ZN (new_n7912_),
	   .A2 (net_6568),
	   .A1 (new_n6973_) );
   NAND2_X1 g1181 (
	   .ZN (new_n7911_1_),
	   .A2 (new_n6980_),
	   .A1 (new_n7910_) );
   NAND4_X1 g1180 (
	   .ZN (new_n7910_),
	   .A4 (new_n7909_),
	   .A3 (new_n7908_),
	   .A2 (new_n7907_),
	   .A1 (new_n7906_1_) );
   NAND3_X1 g1179 (
	   .ZN (new_n7909_),
	   .A3 (_net_6689),
	   .A2 (net_6666),
	   .A1 (_net_6688) );
   NAND3_X1 g1178 (
	   .ZN (new_n7908_),
	   .A3 (net_6634),
	   .A2 (_net_6689),
	   .A1 (new_n7004_) );
   NAND3_X1 g1177 (
	   .ZN (new_n7907_),
	   .A3 (_net_6688),
	   .A2 (net_6602),
	   .A1 (new_n7002_) );
   NAND2_X1 g1176 (
	   .ZN (new_n7906_1_),
	   .A2 (net_6570),
	   .A1 (new_n6973_) );
   AND3_X1 g1175 (
	   .ZN (new_n7905_),
	   .A3 (new_n7904_),
	   .A2 (new_n7903_),
	   .A1 (new_n7902_1_) );
   NAND4_X1 g1174 (
	   .ZN (new_n7904_),
	   .A4 (new_n6987_),
	   .A3 (_net_6687),
	   .A2 (net_6646),
	   .A1 (new_n7118_) );
   NAND4_X1 g1173 (
	   .ZN (new_n7903_),
	   .A4 (new_n6990_1_),
	   .A3 (net_6582),
	   .A2 (_net_6687),
	   .A1 (new_n7115_) );
   NAND4_X1 g1172 (
	   .ZN (new_n7902_1_),
	   .A4 (new_n6989_),
	   .A3 (net_6614),
	   .A2 (_net_6687),
	   .A1 (new_n7115_) );
   CLKBUF_X1 g1171 (
	   .Z (n1515),
	   .A (net_6619) );
   CLKBUF_X1 g1170 (
	   .Z (n1510),
	   .A (_net_7824) );
   CLKBUF_X1 g1169 (
	   .Z (n1506),
	   .A (net_7550) );
   MUX2_X1 g1168 (
	   .Z (n1501),
	   .S (new_n7285_),
	   .B (_net_7698),
	   .A (_net_7800) );
   AOI21_X1 g1167 (
	   .ZN (n1496),
	   .B2 (net_307),
	   .B1 (_net_6007),
	   .A (new_n7896_) );
   NAND3_X1 g1166 (
	   .ZN (new_n7896_),
	   .A3 (_net_6006),
	   .A2 (new_n7895_),
	   .A1 (new_n7655_) );
   INV_X1 g1165 (
	   .ZN (new_n7895_),
	   .A (net_7754) );
   CLKBUF_X1 g1164 (
	   .Z (n1491),
	   .A (_net_7803) );
   AOI21_X1 g1163 (
	   .ZN (n1487),
	   .B2 (new_n7892_),
	   .B1 (new_n7891_),
	   .A (new_n7428_) );
   INV_X1 g1162 (
	   .ZN (new_n7892_),
	   .A (net_297) );
   INV_X1 g1161 (
	   .ZN (new_n7891_),
	   .A (_net_7746) );
   CLKBUF_X1 g1160 (
	   .Z (n1482),
	   .A (x1417) );
   CLKBUF_X1 g1159 (
	   .Z (n1478),
	   .A (_net_6106) );
   CLKBUF_X1 g1158 (
	   .Z (n1474),
	   .A (net_6612) );
   CLKBUF_X1 g1157 (
	   .Z (n1469),
	   .A (net_6392) );
   CLKBUF_X1 g1156 (
	   .Z (n1465),
	   .A (_net_7821) );
   CLKBUF_X1 g1155 (
	   .Z (n1460),
	   .A (_net_6132) );
   CLKBUF_X1 g1154 (
	   .Z (n1455),
	   .A (_net_7803) );
   MUX2_X1 g1153 (
	   .Z (n1451),
	   .S (new_n6823_),
	   .B (_net_6044),
	   .A (_net_7806) );
   CLKBUF_X1 g1152 (
	   .Z (n1446),
	   .A (_net_7813) );
   MUX2_X1 g1151 (
	   .Z (n1442),
	   .S (new_n7609_),
	   .B (_net_7565),
	   .A (new_n7523_) );
   CLKBUF_X1 g1150 (
	   .Z (n1438),
	   .A (net_6745) );
   NOR3_X1 g1149 (
	   .ZN (n1433),
	   .A3 (new_n6821_),
	   .A2 (x1322),
	   .A1 (new_n7878_1_) );
   NAND2_X1 g1148 (
	   .ZN (new_n7878_1_),
	   .A2 (x1261),
	   .A1 (new_n6819_) );
   OAI21_X1 g1147 (
	   .ZN (n1428),
	   .B2 (new_n7736_),
	   .B1 (new_n7876_),
	   .A (new_n7875_1_) );
   INV_X1 g1146 (
	   .ZN (new_n7876_),
	   .A (_net_7497) );
   NAND2_X1 g1145 (
	   .ZN (new_n7875_1_),
	   .A2 (new_n7874_),
	   .A1 (new_n7733_) );
   OAI21_X1 g1144 (
	   .ZN (new_n7874_),
	   .B2 (new_n7873_),
	   .B1 (new_n7034_),
	   .A (new_n7872_) );
   INV_X1 g1143 (
	   .ZN (new_n7873_),
	   .A (net_7385) );
   AOI22_X1 g1142 (
	   .ZN (new_n7872_),
	   .B2 (_net_281),
	   .B1 (net_346),
	   .A2 (net_348),
	   .A1 (_net_280) );
   CLKBUF_X1 g1141 (
	   .Z (n1423),
	   .A (_net_7809) );
   OAI21_X1 g1140 (
	   .ZN (n1419),
	   .B2 (new_n6957_1_),
	   .B1 (new_n7869_),
	   .A (new_n7868_) );
   INV_X1 g1139 (
	   .ZN (new_n7869_),
	   .A (_net_7253) );
   NAND2_X1 g1138 (
	   .ZN (new_n7868_),
	   .A2 (new_n7255_),
	   .A1 (new_n6949_) );
   CLKBUF_X1 g1137 (
	   .Z (n1414),
	   .A (_net_7815) );
   AOI21_X1 g1136 (
	   .ZN (n1410),
	   .B2 (new_n7865_),
	   .B1 (new_n7862_),
	   .A (new_n7855_) );
   OAI211_X1 g1135 (
	   .ZN (new_n7865_),
	   .C2 (new_n7859_),
	   .C1 (new_n7858_1_),
	   .B (new_n7864_),
	   .A (new_n7863_1_) );
   INV_X1 g1134 (
	   .ZN (new_n7864_),
	   .A (new_n7861_) );
   INV_X1 g1133 (
	   .ZN (new_n7863_1_),
	   .A (_net_6558) );
   OAI21_X1 g1132 (
	   .ZN (new_n7862_),
	   .B2 (new_n7861_),
	   .B1 (new_n7860_),
	   .A (_net_6558) );
   NOR2_X1 g1131 (
	   .ZN (new_n7861_),
	   .A2 (_net_6552),
	   .A1 (new_n7857_) );
   NOR2_X1 g1130 (
	   .ZN (new_n7860_),
	   .A2 (new_n7859_),
	   .A1 (new_n7858_1_) );
   INV_X1 g1129 (
	   .ZN (new_n7859_),
	   .A (_net_6552) );
   XNOR2_X1 g1128 (
	   .ZN (new_n7858_1_),
	   .B (new_n7857_),
	   .A (new_n7856_) );
   INV_X1 g1127 (
	   .ZN (new_n7857_),
	   .A (_net_6555) );
   NAND2_X1 g1126 (
	   .ZN (new_n7856_),
	   .A2 (_net_6554),
	   .A1 (_net_6553) );
   NAND4_X1 g1125 (
	   .ZN (new_n7855_),
	   .A4 (new_n7854_),
	   .A3 (new_n7853_1_),
	   .A2 (new_n7851_),
	   .A1 (new_n7848_1_) );
   OAI21_X1 g1124 (
	   .ZN (new_n7854_),
	   .B2 (new_n6761_1_),
	   .B1 (n8472),
	   .A (_net_6552) );
   OR2_X1 g1123 (
	   .ZN (new_n7853_1_),
	   .A2 (_net_6552),
	   .A1 (n8472) );
   XNOR2_X1 g1122 (
	   .ZN (n8472),
	   .B (_net_6553),
	   .A (net_6556) );
   NAND2_X1 g1121 (
	   .ZN (new_n7851_),
	   .A2 (new_n7850_),
	   .A1 (new_n7849_) );
   INV_X1 g1120 (
	   .ZN (new_n7850_),
	   .A (_net_6557) );
   XNOR2_X1 g1119 (
	   .ZN (new_n7849_),
	   .B (_net_6554),
	   .A (new_n6778_) );
   NAND2_X1 g1118 (
	   .ZN (new_n7848_1_),
	   .A2 (_net_6557),
	   .A1 (new_n7847_) );
   XNOR2_X1 g1117 (
	   .ZN (new_n7847_),
	   .B (new_n6787_),
	   .A (new_n6778_) );
   NAND3_X1 g1116 (
	   .ZN (n1405),
	   .A3 (new_n7845_1_),
	   .A2 (new_n7835_1_),
	   .A1 (new_n7818_1_) );
   AOI22_X1 g1115 (
	   .ZN (new_n7845_1_),
	   .B2 (net_7225),
	   .B1 (new_n7844_),
	   .A2 (new_n7842_),
	   .A1 (new_n7837_) );
   NOR3_X2 g1114 (
	   .ZN (new_n7844_),
	   .A3 (new_n7843_),
	   .A2 (new_n7811_),
	   .A1 (new_n7687_) );
   NAND3_X1 g1113 (
	   .ZN (new_n7843_),
	   .A3 (_net_7228),
	   .A2 (_net_7227),
	   .A1 (_net_7229) );
   NAND4_X1 g1112 (
	   .ZN (new_n7842_),
	   .A4 (new_n7841_),
	   .A3 (new_n7840_1_),
	   .A2 (new_n7839_),
	   .A1 (new_n7838_) );
   NAND3_X1 g1111 (
	   .ZN (new_n7841_),
	   .A3 (_net_7228),
	   .A2 (net_7209),
	   .A1 (_net_7229) );
   NAND3_X1 g1110 (
	   .ZN (new_n7840_1_),
	   .A3 (net_7177),
	   .A2 (_net_7229),
	   .A1 (new_n7823_) );
   NAND3_X1 g1109 (
	   .ZN (new_n7839_),
	   .A3 (_net_7228),
	   .A2 (net_7145),
	   .A1 (new_n7821_) );
   NAND2_X1 g1108 (
	   .ZN (new_n7838_),
	   .A2 (net_7113),
	   .A1 (new_n7819_) );
   BUF_X4 g1107 (
	   .Z (new_n7837_),
	   .A (new_n7836_) );
   NOR3_X1 g1106 (
	   .ZN (new_n7836_),
	   .A3 (_net_7227),
	   .A2 (new_n7811_),
	   .A1 (new_n7687_) );
   AND3_X1 g1105 (
	   .ZN (new_n7835_1_),
	   .A3 (new_n7834_),
	   .A2 (new_n7833_),
	   .A1 (new_n7827_) );
   NAND2_X1 g1104 (
	   .ZN (new_n7834_),
	   .A2 (_net_6182),
	   .A1 (new_n7694_) );
   NAND2_X1 g1103 (
	   .ZN (new_n7833_),
	   .A2 (new_n7689_),
	   .A1 (new_n7832_) );
   NAND4_X1 g1102 (
	   .ZN (new_n7832_),
	   .A4 (new_n7831_1_),
	   .A3 (new_n7830_),
	   .A2 (new_n7829_),
	   .A1 (new_n7828_) );
   NAND3_X1 g1101 (
	   .ZN (new_n7831_1_),
	   .A3 (_net_7228),
	   .A2 (net_7213),
	   .A1 (_net_7229) );
   NAND3_X1 g1100 (
	   .ZN (new_n7830_),
	   .A3 (net_7181),
	   .A2 (_net_7229),
	   .A1 (new_n7823_) );
   NAND3_X1 g1099 (
	   .ZN (new_n7829_),
	   .A3 (_net_7228),
	   .A2 (net_7149),
	   .A1 (new_n7821_) );
   NAND2_X1 g1098 (
	   .ZN (new_n7828_),
	   .A2 (net_7117),
	   .A1 (new_n7819_) );
   NAND2_X1 g1097 (
	   .ZN (new_n7827_),
	   .A2 (new_n7701_),
	   .A1 (new_n7826_1_) );
   NAND4_X1 g1096 (
	   .ZN (new_n7826_1_),
	   .A4 (new_n7825_),
	   .A3 (new_n7824_),
	   .A2 (new_n7822_1_),
	   .A1 (new_n7820_) );
   NAND3_X1 g1095 (
	   .ZN (new_n7825_),
	   .A3 (_net_7228),
	   .A2 (net_7211),
	   .A1 (_net_7229) );
   NAND3_X1 g1094 (
	   .ZN (new_n7824_),
	   .A3 (_net_7229),
	   .A2 (net_7179),
	   .A1 (new_n7823_) );
   BUF_X4 g1093 (
	   .Z (new_n7823_),
	   .A (new_n7675_) );
   NAND3_X1 g1092 (
	   .ZN (new_n7822_1_),
	   .A3 (_net_7228),
	   .A2 (net_7147),
	   .A1 (new_n7821_) );
   BUF_X4 g1091 (
	   .Z (new_n7821_),
	   .A (new_n7674_) );
   NAND2_X1 g1090 (
	   .ZN (new_n7820_),
	   .A2 (net_7115),
	   .A1 (new_n7819_) );
   BUF_X4 g1089 (
	   .Z (new_n7819_),
	   .A (new_n7682_) );
   AND3_X1 g1088 (
	   .ZN (new_n7818_1_),
	   .A3 (new_n7817_),
	   .A2 (new_n7815_1_),
	   .A1 (new_n7814_) );
   NAND4_X1 g1087 (
	   .ZN (new_n7817_),
	   .A4 (new_n7678_),
	   .A3 (net_7193),
	   .A2 (_net_7227),
	   .A1 (new_n7816_) );
   BUF_X4 g1086 (
	   .Z (new_n7816_),
	   .A (new_n7812_) );
   NAND4_X1 g1085 (
	   .ZN (new_n7815_1_),
	   .A4 (new_n7683_),
	   .A3 (net_7129),
	   .A2 (_net_7227),
	   .A1 (new_n7813_) );
   NAND4_X1 g1084 (
	   .ZN (new_n7814_),
	   .A4 (new_n7681_1_),
	   .A3 (net_7161),
	   .A2 (_net_7227),
	   .A1 (new_n7813_) );
   BUF_X4 g1083 (
	   .Z (new_n7813_),
	   .A (new_n7812_) );
   NOR2_X2 g1082 (
	   .ZN (new_n7812_),
	   .A2 (new_n7811_),
	   .A1 (new_n7687_) );
   INV_X1 g1081 (
	   .ZN (new_n7811_),
	   .A (new_n7810_1_) );
   NOR2_X1 g1080 (
	   .ZN (new_n7810_1_),
	   .A2 (_net_6041),
	   .A1 (_net_6042) );
   CLKBUF_X1 g1079 (
	   .Z (n1400),
	   .A (_net_7794) );
   AND2_X1 g1078 (
	   .ZN (n1396),
	   .A2 (_net_6189),
	   .A1 (new_n7239_) );
   MUX2_X1 g1077 (
	   .Z (n1391),
	   .S (new_n7545_),
	   .B (_net_7658),
	   .A (new_n7806_1_) );
   OAI21_X1 g1076 (
	   .ZN (new_n7806_1_),
	   .B2 (new_n7805_),
	   .B1 (new_n7020_),
	   .A (new_n7804_) );
   INV_X1 g1075 (
	   .ZN (new_n7805_),
	   .A (net_7546) );
   AOI22_X1 g1074 (
	   .ZN (new_n7804_),
	   .B2 (_net_291),
	   .B1 (net_378),
	   .A2 (_net_292),
	   .A1 (net_376) );
   CLKBUF_X1 g1073 (
	   .Z (n1386),
	   .A (net_6400) );
   CLKBUF_X1 g1072 (
	   .Z (n1383),
	   .A (net_6694) );
   CLKBUF_X1 g1071 (
	   .Z (n1378),
	   .A (_net_5960) );
   MUX2_X1 g1070 (
	   .Z (n1373),
	   .S (new_n7437_1_),
	   .B (_net_5997),
	   .A (_net_7803) );
   AOI21_X1 g1069 (
	   .ZN (n1368),
	   .B2 (new_n7798_1_),
	   .B1 (new_n7797_),
	   .A (new_n6867_1_) );
   AOI21_X1 g1068 (
	   .ZN (new_n7798_1_),
	   .B2 (new_n7796_),
	   .B1 (new_n7795_),
	   .A (_net_5972) );
   OAI21_X1 g1067 (
	   .ZN (new_n7797_),
	   .B2 (new_n7796_),
	   .B1 (new_n7795_),
	   .A (new_n7794_) );
   INV_X1 g1066 (
	   .ZN (new_n7796_),
	   .A (_net_5974) );
   NOR2_X1 g1065 (
	   .ZN (new_n7795_),
	   .A2 (_net_5973),
	   .A1 (_net_6021) );
   INV_X1 g1064 (
	   .ZN (new_n7794_),
	   .A (_net_6022) );
   NAND2_X1 g1063 (
	   .ZN (n1363),
	   .A2 (new_n7792_),
	   .A1 (new_n7791_) );
   AOI22_X1 g1062 (
	   .ZN (new_n7792_),
	   .B2 (net_7517),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7485) );
   AOI22_X1 g1061 (
	   .ZN (new_n7791_),
	   .B2 (_net_7421),
	   .B1 (new_n7298_),
	   .A2 (net_7453),
	   .A1 (new_n7296_) );
   CLKBUF_X1 g1060 (
	   .Z (n1359),
	   .A (net_7234) );
   CLKBUF_X1 g1059 (
	   .Z (n1355),
	   .A (net_6877) );
   AND2_X1 g1058 (
	   .ZN (n1345),
	   .A2 (_net_6017),
	   .A1 (_net_5975) );
   MUX2_X1 g1057 (
	   .Z (n1340),
	   .S (new_n7285_),
	   .B (_net_7707),
	   .A (_net_7809) );
   MUX2_X1 g1056 (
	   .Z (n1335),
	   .S (new_n7437_1_),
	   .B (_net_5991),
	   .A (_net_7800) );
   CLKBUF_X1 g1055 (
	   .Z (n1331),
	   .A (net_6859) );
   CLKBUF_X1 g1054 (
	   .Z (n1326),
	   .A (_net_7820) );
   CLKBUF_X1 g1053 (
	   .Z (n1322),
	   .A (_net_7798) );
   CLKBUF_X1 g1052 (
	   .Z (n1318),
	   .A (_net_7812) );
   MUX2_X1 g1051 (
	   .Z (n1314),
	   .S (new_n7437_1_),
	   .B (_net_6000),
	   .A (_net_7806) );
   XNOR2_X1 g1050 (
	   .ZN (n1309),
	   .B (new_n7227_),
	   .A (new_n7779_1_) );
   XNOR2_X1 g1049 (
	   .ZN (new_n7779_1_),
	   .B (_net_6692),
	   .A (_net_6689) );
   CLKBUF_X1 g1048 (
	   .Z (n1305),
	   .A (net_7395) );
   CLKBUF_X1 g1047 (
	   .Z (n1300),
	   .A (_net_7803) );
   OAI21_X1 g1046 (
	   .ZN (n1295),
	   .B2 (new_n7225_),
	   .B1 (new_n7775_),
	   .A (new_n7774_) );
   INV_X1 g1045 (
	   .ZN (new_n7775_),
	   .A (_net_7315) );
   NAND2_X1 g1044 (
	   .ZN (new_n7774_),
	   .A2 (new_n7773_1_),
	   .A1 (new_n7222_) );
   OAI21_X1 g1043 (
	   .ZN (new_n7773_1_),
	   .B2 (new_n7772_),
	   .B1 (new_n6952_1_),
	   .A (new_n7771_) );
   INV_X1 g1042 (
	   .ZN (new_n7772_),
	   .A (net_7235) );
   AOI22_X1 g1041 (
	   .ZN (new_n7771_),
	   .B2 (net_327),
	   .B1 (_net_270),
	   .A2 (_net_269),
	   .A1 (net_329) );
   CLKBUF_X1 g1040 (
	   .Z (n1291),
	   .A (net_6574) );
   CLKBUF_X1 g1039 (
	   .Z (n1287),
	   .A (net_7119) );
   OAI21_X1 g1038 (
	   .ZN (n1282),
	   .B2 (new_n7767_),
	   .B1 (new_n7024_),
	   .A (new_n7766_) );
   INV_X1 g1037 (
	   .ZN (new_n7767_),
	   .A (_net_263) );
   INV_X1 g1036 (
	   .ZN (new_n7766_),
	   .A (_net_299) );
   NOR2_X1 g1035 (
	   .ZN (n1277),
	   .A2 (new_n7275_1_),
	   .A1 (new_n7035_) );
   MUX2_X1 g1034 (
	   .Z (n1272),
	   .S (new_n7538_),
	   .B (_net_273),
	   .A (net_7799) );
   MUX2_X1 g1033 (
	   .Z (n1267),
	   .S (new_n7029_),
	   .B (_net_7590),
	   .A (new_n7762_) );
   OAI21_X1 g1032 (
	   .ZN (new_n7762_),
	   .B2 (new_n7761_),
	   .B1 (new_n7020_),
	   .A (new_n7760_1_) );
   INV_X1 g1031 (
	   .ZN (new_n7761_),
	   .A (net_7542) );
   AOI22_X1 g1030 (
	   .ZN (new_n7760_1_),
	   .B2 (net_374),
	   .B1 (_net_291),
	   .A2 (_net_292),
	   .A1 (net_372) );
   CLKBUF_X1 g1029 (
	   .Z (n1262),
	   .A (_net_6158) );
   CLKBUF_X1 g1028 (
	   .Z (n1258),
	   .A (net_7019) );
   OAI21_X1 g1027 (
	   .ZN (n1253),
	   .B2 (new_n7736_),
	   .B1 (new_n7756_1_),
	   .A (new_n7755_) );
   INV_X1 g1026 (
	   .ZN (new_n7756_1_),
	   .A (_net_7512) );
   NAND2_X1 g1025 (
	   .ZN (new_n7755_),
	   .A2 (new_n7754_),
	   .A1 (new_n7733_) );
   OAI21_X1 g1024 (
	   .ZN (new_n7754_),
	   .B2 (new_n7753_),
	   .B1 (new_n7034_),
	   .A (new_n7752_) );
   INV_X1 g1023 (
	   .ZN (new_n7753_),
	   .A (net_7400) );
   AOI22_X1 g1022 (
	   .ZN (new_n7752_),
	   .B2 (_net_280),
	   .B1 (net_363),
	   .A2 (_net_281),
	   .A1 (net_361) );
   CLKBUF_X1 g1021 (
	   .Z (n1248),
	   .A (_net_7794) );
   CLKBUF_X1 g1020 (
	   .Z (n1244),
	   .A (net_6395) );
   CLKBUF_X1 g1019 (
	   .Z (n1240),
	   .A (_net_7820) );
   AND2_X1 g1018 (
	   .ZN (n1236),
	   .A2 (net_381),
	   .A1 (new_n7747_) );
   BUF_X2 g1017 (
	   .Z (new_n7747_),
	   .A (new_n7262_) );
   CLKBUF_X1 g1016 (
	   .Z (n1232),
	   .A (_net_7795) );
   AOI21_X1 g1015 (
	   .ZN (n1228),
	   .B2 (new_n7744_),
	   .B1 (new_n7376_1_),
	   .A (new_n7428_) );
   INV_X1 g1014 (
	   .ZN (new_n7744_),
	   .A (_net_6016) );
   CLKBUF_X1 g1013 (
	   .Z (n1224),
	   .A (net_6608) );
   AOI21_X1 g1012 (
	   .ZN (n1219),
	   .B2 (new_n7739_),
	   .B1 (new_n7741_1_),
	   .A (new_n7740_) );
   INV_X1 g1011 (
	   .ZN (new_n7741_1_),
	   .A (_net_7428) );
   NOR2_X1 g1010 (
	   .ZN (new_n7740_),
	   .A2 (n595),
	   .A1 (new_n7739_) );
   BUF_X4 g1009 (
	   .Z (new_n7739_),
	   .A (new_n7738_) );
   NAND2_X2 g1008 (
	   .ZN (new_n7738_),
	   .A2 (new_n7643_),
	   .A1 (new_n6892_) );
   OAI21_X1 g1007 (
	   .ZN (n1214),
	   .B2 (new_n7736_),
	   .B1 (new_n7735_),
	   .A (new_n7734_) );
   BUF_X4 g1006 (
	   .Z (new_n7736_),
	   .A (new_n7732_1_) );
   INV_X1 g1005 (
	   .ZN (new_n7735_),
	   .A (_net_7503) );
   NAND2_X1 g1004 (
	   .ZN (new_n7734_),
	   .A2 (new_n7484_),
	   .A1 (new_n7733_) );
   BUF_X4 g1003 (
	   .Z (new_n7733_),
	   .A (new_n7732_1_) );
   BUF_X4 g1002 (
	   .Z (new_n7732_1_),
	   .A (new_n7731_) );
   AND2_X1 g1001 (
	   .ZN (new_n7731_),
	   .A2 (new_n7730_),
	   .A1 (new_n6892_) );
   NOR2_X1 g1000 (
	   .ZN (new_n7730_),
	   .A2 (new_n7268_),
	   .A1 (new_n6893_) );
   CLKBUF_X1 g0999 (
	   .Z (n1210),
	   .A (net_6845) );
   CLKBUF_X1 g0998 (
	   .Z (n1205),
	   .A (_net_7814) );
   CLKBUF_X1 g0997 (
	   .Z (n1200),
	   .A (_net_6064) );
   CLKBUF_X1 g0996 (
	   .Z (n1195),
	   .A (_net_7822) );
   CLKBUF_X1 g0995 (
	   .Z (n1191),
	   .A (_net_7823) );
   CLKBUF_X1 g0994 (
	   .Z (n1187),
	   .A (net_6400) );
   CLKBUF_X1 g0993 (
	   .Z (n1183),
	   .A (net_144) );
   NAND3_X1 g0992 (
	   .ZN (n1178),
	   .A3 (new_n7721_),
	   .A2 (new_n7720_),
	   .A1 (new_n7711_) );
   AOI22_X1 g0991 (
	   .ZN (new_n7721_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6948),
	   .A2 (new_n6860_1_),
	   .A1 (new_n6879_) );
   AND3_X1 g0990 (
	   .ZN (new_n7720_),
	   .A3 (new_n7719_1_),
	   .A2 (new_n7718_),
	   .A1 (new_n7717_) );
   NAND2_X1 g0989 (
	   .ZN (new_n7719_1_),
	   .A2 (_net_6135),
	   .A1 (new_n6869_) );
   NAND2_X1 g0988 (
	   .ZN (new_n7718_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n6851_) );
   NAND2_X1 g0987 (
	   .ZN (new_n7717_),
	   .A2 (new_n6854_),
	   .A1 (new_n7716_) );
   NAND4_X1 g0986 (
	   .ZN (new_n7716_),
	   .A4 (new_n7715_),
	   .A3 (new_n7714_1_),
	   .A2 (new_n7713_),
	   .A1 (new_n7712_) );
   NAND3_X1 g0985 (
	   .ZN (new_n7715_),
	   .A3 (net_6936),
	   .A2 (_net_6958),
	   .A1 (_net_6959) );
   NAND3_X1 g0984 (
	   .ZN (new_n7714_1_),
	   .A3 (_net_6959),
	   .A2 (net_6904),
	   .A1 (new_n6848_) );
   NAND3_X1 g0983 (
	   .ZN (new_n7713_),
	   .A3 (_net_6958),
	   .A2 (net_6872),
	   .A1 (new_n6846_) );
   NAND2_X1 g0982 (
	   .ZN (new_n7712_),
	   .A2 (net_6840),
	   .A1 (new_n6844_) );
   AND3_X1 g0981 (
	   .ZN (new_n7711_),
	   .A3 (new_n7710_),
	   .A2 (new_n7709_1_),
	   .A1 (new_n7708_) );
   NAND4_X1 g0980 (
	   .ZN (new_n7710_),
	   .A4 (new_n6841_),
	   .A3 (net_6916),
	   .A2 (_net_6957),
	   .A1 (new_n6838_) );
   NAND4_X1 g0979 (
	   .ZN (new_n7709_1_),
	   .A4 (new_n6836_1_),
	   .A3 (_net_6957),
	   .A2 (net_6852),
	   .A1 (new_n6830_) );
   NAND4_X1 g0978 (
	   .ZN (new_n7708_),
	   .A4 (new_n6833_),
	   .A3 (net_6884),
	   .A2 (_net_6957),
	   .A1 (new_n6830_) );
   NOR2_X1 g0977 (
	   .ZN (n1173),
	   .A2 (new_n7594_),
	   .A1 (new_n7035_) );
   CLKBUF_X1 g0976 (
	   .Z (n1168),
	   .A (net_6398) );
   AND2_X1 g0975 (
	   .ZN (n1163),
	   .A2 (net_381),
	   .A1 (new_n7262_) );
   CLKBUF_X1 g0974 (
	   .Z (n1158),
	   .A (_net_6066) );
   NAND2_X1 g0973 (
	   .ZN (n1153),
	   .A2 (new_n7702_),
	   .A1 (new_n7695_1_) );
   NAND2_X1 g0972 (
	   .ZN (new_n7702_),
	   .A2 (new_n7701_),
	   .A1 (new_n7698_) );
   BUF_X4 g0971 (
	   .Z (new_n7701_),
	   .A (new_n7700_1_) );
   NOR2_X1 g0970 (
	   .ZN (new_n7700_1_),
	   .A2 (new_n7699_),
	   .A1 (new_n7687_) );
   INV_X1 g0969 (
	   .ZN (new_n7699_),
	   .A (_net_6041) );
   NAND2_X1 g0968 (
	   .ZN (new_n7698_),
	   .A2 (new_n7697_),
	   .A1 (new_n7696_) );
   AOI22_X1 g0967 (
	   .ZN (new_n7697_),
	   .B2 (net_7100),
	   .B1 (new_n7683_),
	   .A2 (net_7132),
	   .A1 (new_n7681_1_) );
   AOI22_X1 g0966 (
	   .ZN (new_n7696_),
	   .B2 (net_7164),
	   .B1 (new_n7678_),
	   .A2 (new_n7676_1_),
	   .A1 (net_7196) );
   AOI22_X1 g0965 (
	   .ZN (new_n7695_1_),
	   .B2 (new_n7694_),
	   .B1 (_net_6167),
	   .A2 (new_n7690_),
	   .A1 (new_n7685_) );
   BUF_X4 g0964 (
	   .Z (new_n7694_),
	   .A (new_n7693_) );
   INV_X1 g0963 (
	   .ZN (new_n7693_),
	   .A (new_n7692_) );
   NAND2_X1 g0962 (
	   .ZN (new_n7692_),
	   .A2 (_net_6039),
	   .A1 (new_n7691_1_) );
   NAND3_X1 g0961 (
	   .ZN (new_n7691_1_),
	   .A3 (net_6056),
	   .A2 (_net_7791),
	   .A1 (new_n7686_1_) );
   BUF_X4 g0960 (
	   .Z (new_n7690_),
	   .A (new_n7689_) );
   NOR2_X1 g0959 (
	   .ZN (new_n7689_),
	   .A2 (new_n7688_),
	   .A1 (new_n7687_) );
   INV_X1 g0958 (
	   .ZN (new_n7688_),
	   .A (_net_6042) );
   NAND4_X1 g0957 (
	   .ZN (new_n7687_),
	   .A4 (_net_6039),
	   .A3 (net_6056),
	   .A2 (_net_7791),
	   .A1 (new_n7686_1_) );
   INV_X1 g0956 (
	   .ZN (new_n7686_1_),
	   .A (_net_7759) );
   NAND2_X1 g0955 (
	   .ZN (new_n7685_),
	   .A2 (new_n7684_),
	   .A1 (new_n7679_) );
   AOI22_X1 g0954 (
	   .ZN (new_n7684_),
	   .B2 (net_7102),
	   .B1 (new_n7683_),
	   .A2 (net_7134),
	   .A1 (new_n7681_1_) );
   BUF_X4 g0953 (
	   .Z (new_n7683_),
	   .A (new_n7682_) );
   NOR2_X1 g0952 (
	   .ZN (new_n7682_),
	   .A2 (_net_7228),
	   .A1 (_net_7229) );
   BUF_X4 g0951 (
	   .Z (new_n7681_1_),
	   .A (new_n7680_) );
   NOR2_X1 g0950 (
	   .ZN (new_n7680_),
	   .A2 (_net_7229),
	   .A1 (new_n7675_) );
   AOI22_X1 g0949 (
	   .ZN (new_n7679_),
	   .B2 (net_7166),
	   .B1 (new_n7678_),
	   .A2 (new_n7676_1_),
	   .A1 (net_7198) );
   BUF_X4 g0948 (
	   .Z (new_n7678_),
	   .A (new_n7677_) );
   NOR2_X1 g0947 (
	   .ZN (new_n7677_),
	   .A2 (_net_7228),
	   .A1 (new_n7674_) );
   NOR2_X1 g0946 (
	   .ZN (new_n7676_1_),
	   .A2 (new_n7675_),
	   .A1 (new_n7674_) );
   INV_X1 g0945 (
	   .ZN (new_n7675_),
	   .A (_net_7228) );
   INV_X1 g0944 (
	   .ZN (new_n7674_),
	   .A (_net_7229) );
   CLKBUF_X1 g0943 (
	   .Z (n1148),
	   .A (_net_7815) );
   CLKBUF_X1 g0942 (
	   .Z (n1144),
	   .A (_net_6099) );
   CLKBUF_X1 g0941 (
	   .Z (n1140),
	   .A (net_6986) );
   OAI21_X1 g0940 (
	   .ZN (n1135),
	   .B2 (new_n7258_),
	   .B1 (new_n7669_),
	   .A (new_n7668_) );
   INV_X1 g0939 (
	   .ZN (new_n7669_),
	   .A (_net_7299) );
   NAND2_X1 g0938 (
	   .ZN (new_n7668_),
	   .A2 (new_n7667_),
	   .A1 (new_n7252_1_) );
   OAI21_X1 g0937 (
	   .ZN (new_n7667_),
	   .B2 (new_n7666_1_),
	   .B1 (new_n6952_1_),
	   .A (new_n7665_) );
   INV_X1 g0936 (
	   .ZN (new_n7666_1_),
	   .A (net_331) );
   AOI22_X1 g0935 (
	   .ZN (new_n7665_),
	   .B2 (net_343),
	   .B1 (_net_270),
	   .A2 (_net_269),
	   .A1 (net_345) );
   CLKBUF_X1 g0934 (
	   .Z (n1130),
	   .A (_net_7809) );
   AOI21_X1 g0933 (
	   .ZN (n1125),
	   .B2 (new_n7326_1_),
	   .B1 (new_n7662_),
	   .A (new_n7661_1_) );
   INV_X1 g0932 (
	   .ZN (new_n7662_),
	   .A (_net_7274) );
   NOR2_X1 g0931 (
	   .ZN (new_n7661_1_),
	   .A2 (n4263),
	   .A1 (new_n7326_1_) );
   AND2_X1 g0930 (
	   .ZN (n4263),
	   .A2 (net_338),
	   .A1 (new_n7102_1_) );
   CLKBUF_X1 g0929 (
	   .Z (n1121),
	   .A (net_6847) );
   AOI21_X1 g0928 (
	   .ZN (n1116),
	   .B2 (net_308),
	   .B1 (_net_5996),
	   .A (new_n7657_) );
   NAND3_X1 g0927 (
	   .ZN (new_n7657_),
	   .A3 (_net_5995),
	   .A2 (new_n7656_),
	   .A1 (new_n7655_) );
   INV_X1 g0926 (
	   .ZN (new_n7656_),
	   .A (net_7752) );
   AND2_X2 g0925 (
	   .ZN (new_n7655_),
	   .A2 (_net_7791),
	   .A1 (net_303) );
   CLKBUF_X1 g0924 (
	   .Z (n1111),
	   .A (_net_6183) );
   OAI21_X1 g0923 (
	   .ZN (n1106),
	   .B2 (new_n7652_),
	   .B1 (new_n7651_),
	   .A (new_n7650_) );
   BUF_X4 g0922 (
	   .Z (new_n7652_),
	   .A (new_n7645_) );
   INV_X1 g0921 (
	   .ZN (new_n7651_),
	   .A (_net_7412) );
   NAND2_X1 g0920 (
	   .ZN (new_n7650_),
	   .A2 (new_n7649_1_),
	   .A1 (new_n7646_) );
   OAI221_X1 g0919 (
	   .ZN (new_n7649_1_),
	   .C2 (new_n7648_),
	   .C1 (new_n6902_1_),
	   .B2 (new_n6901_),
	   .B1 (new_n6933_),
	   .A (new_n7647_) );
   INV_X1 g0918 (
	   .ZN (new_n7648_),
	   .A (net_359) );
   NAND2_X1 g0917 (
	   .ZN (new_n7647_),
	   .A2 (net_7396),
	   .A1 (new_n6898_) );
   BUF_X4 g0916 (
	   .Z (new_n7646_),
	   .A (new_n7645_) );
   BUF_X4 g0915 (
	   .Z (new_n7645_),
	   .A (new_n7644_1_) );
   AND2_X1 g0914 (
	   .ZN (new_n7644_1_),
	   .A2 (new_n7643_),
	   .A1 (new_n6892_) );
   NOR2_X1 g0913 (
	   .ZN (new_n7643_),
	   .A2 (_net_7533),
	   .A1 (_net_7534) );
   CLKBUF_X1 g0912 (
	   .Z (n1102),
	   .A (net_6856) );
   CLKBUF_X1 g0911 (
	   .Z (n1097),
	   .A (_net_7801) );
   CLKBUF_X1 g0910 (
	   .Z (n1093),
	   .A (net_6977) );
   CLKBUF_X1 g0909 (
	   .Z (n1089),
	   .A (net_6832) );
   CLKBUF_X1 g0908 (
	   .Z (n1085),
	   .A (net_6461) );
   CLKBUF_X1 g0907 (
	   .Z (n1081),
	   .A (net_7010) );
   CLKBUF_X1 g0906 (
	   .Z (n1077),
	   .A (net_7004) );
   AND2_X1 g0905 (
	   .ZN (n1072),
	   .A2 (_net_6285),
	   .A1 (new_n7239_) );
   AOI21_X1 g0904 (
	   .ZN (n1067),
	   .B2 (new_n7633_),
	   .B1 (new_n7632_),
	   .A (new_n6811_) );
   AOI21_X1 g0903 (
	   .ZN (new_n7633_),
	   .B2 (new_n7631_1_),
	   .B1 (new_n7630_),
	   .A (_net_5960) );
   OAI21_X1 g0902 (
	   .ZN (new_n7632_),
	   .B2 (new_n7631_1_),
	   .B1 (new_n7630_),
	   .A (new_n7629_) );
   INV_X1 g0901 (
	   .ZN (new_n7631_1_),
	   .A (_net_5962) );
   NOR2_X1 g0900 (
	   .ZN (new_n7630_),
	   .A2 (_net_5961),
	   .A1 (_net_5988) );
   INV_X1 g0899 (
	   .ZN (new_n7629_),
	   .A (_net_5989) );
   CLKBUF_X1 g0898 (
	   .Z (n1062),
	   .A (_net_7812) );
   NAND3_X1 g0897 (
	   .ZN (n1058),
	   .A3 (new_n7626_1_),
	   .A2 (new_n7625_),
	   .A1 (new_n7616_) );
   NAND4_X1 g0896 (
	   .ZN (new_n7626_1_),
	   .A4 (_net_7697),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   NOR3_X1 g0895 (
	   .ZN (new_n7625_),
	   .A3 (new_n7624_),
	   .A2 (new_n7620_),
	   .A1 (new_n7617_) );
   NAND3_X1 g0894 (
	   .ZN (new_n7624_),
	   .A3 (new_n7623_),
	   .A2 (new_n7622_1_),
	   .A1 (new_n7621_) );
   NAND4_X1 g0893 (
	   .ZN (new_n7623_),
	   .A4 (net_162),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   NAND3_X1 g0892 (
	   .ZN (new_n7622_1_),
	   .A3 (net_199),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   NAND3_X1 g0891 (
	   .ZN (new_n7621_),
	   .A3 (net_236),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   OAI22_X1 g0890 (
	   .ZN (new_n7620_),
	   .B2 (new_n7378_),
	   .B1 (new_n7619_),
	   .A2 (new_n7618_1_),
	   .A1 (new_n7374_) );
   INV_X1 g0889 (
	   .ZN (new_n7619_),
	   .A (_net_7726) );
   INV_X1 g0888 (
	   .ZN (new_n7618_1_),
	   .A (_net_120) );
   AND4_X1 g0887 (
	   .ZN (new_n7617_),
	   .A4 (new_n7371_),
	   .A3 (new_n7360_),
	   .A2 (new_n7369_),
	   .A1 (_net_6034) );
   NOR2_X1 g0886 (
	   .ZN (new_n7616_),
	   .A2 (new_n7615_),
	   .A1 (new_n7613_1_) );
   NOR2_X1 g0885 (
	   .ZN (new_n7615_),
	   .A2 (new_n7614_),
	   .A1 (new_n7366_) );
   INV_X1 g0884 (
	   .ZN (new_n7614_),
	   .A (_net_5990) );
   NOR2_X1 g0883 (
	   .ZN (new_n7613_1_),
	   .A2 (new_n7612_),
	   .A1 (new_n7362_) );
   INV_X1 g0882 (
	   .ZN (new_n7612_),
	   .A (_net_273) );
   CLKBUF_X1 g0881 (
	   .Z (n1053),
	   .A (net_6386) );
   MUX2_X1 g0880 (
	   .Z (n1049),
	   .S (new_n7609_),
	   .B (_net_7578),
	   .A (n3546) );
   BUF_X8 g0879 (
	   .Z (new_n7609_),
	   .A (new_n7608_1_) );
   NAND3_X1 g0878 (
	   .ZN (new_n7608_1_),
	   .A3 (new_n7027_1_),
	   .A2 (new_n7502_),
	   .A1 (new_n7026_) );
   AND2_X1 g0877 (
	   .ZN (n3546),
	   .A2 (net_380),
	   .A1 (new_n7262_) );
   AOI21_X1 g0876 (
	   .ZN (n1044),
	   .B2 (new_n7326_1_),
	   .B1 (new_n7605_),
	   .A (new_n7604_1_) );
   INV_X1 g0875 (
	   .ZN (new_n7605_),
	   .A (_net_7281) );
   NOR2_X1 g0874 (
	   .ZN (new_n7604_1_),
	   .A2 (n6722),
	   .A1 (new_n7326_1_) );
   NOR2_X1 g0873 (
	   .ZN (n6722),
	   .A2 (new_n7602_),
	   .A1 (new_n6952_1_) );
   INV_X1 g0872 (
	   .ZN (new_n7602_),
	   .A (net_345) );
   AND2_X1 g0871 (
	   .ZN (n1039),
	   .A2 (_net_6259),
	   .A1 (new_n7239_) );
   AND2_X1 g0870 (
	   .ZN (n1034),
	   .A2 (net_343),
	   .A1 (new_n7102_1_) );
   NOR2_X1 g0869 (
	   .ZN (n1029),
	   .A2 (new_n7493_),
	   .A1 (new_n6952_1_) );
   OAI21_X1 g0868 (
	   .ZN (n1024),
	   .B2 (new_n7279_),
	   .B1 (new_n7597_),
	   .A (new_n7596_1_) );
   INV_X1 g0867 (
	   .ZN (new_n7597_),
	   .A (_net_7447) );
   NAND2_X1 g0866 (
	   .ZN (new_n7596_1_),
	   .A2 (new_n7595_),
	   .A1 (new_n7272_) );
   OAI221_X1 g0865 (
	   .ZN (new_n7595_),
	   .C2 (new_n6901_),
	   .C1 (new_n7594_),
	   .B2 (new_n6902_1_),
	   .B1 (new_n6900_),
	   .A (new_n7593_) );
   INV_X1 g0864 (
	   .ZN (new_n7594_),
	   .A (net_360) );
   NAND2_X1 g0863 (
	   .ZN (new_n7593_),
	   .A2 (net_7399),
	   .A1 (new_n6898_) );
   CLKBUF_X1 g0862 (
	   .Z (n1020),
	   .A (net_6998) );
   NAND2_X1 g0861 (
	   .ZN (n1015),
	   .A2 (new_n7590_),
	   .A1 (new_n7563_1_) );
   AND4_X1 g0860 (
	   .ZN (new_n7590_),
	   .A4 (new_n7589_),
	   .A3 (new_n7588_),
	   .A2 (new_n7580_),
	   .A1 (new_n7574_) );
   NAND2_X1 g0859 (
	   .ZN (new_n7589_),
	   .A2 (_net_6120),
	   .A1 (new_n7210_) );
   NAND2_X1 g0858 (
	   .ZN (new_n7588_),
	   .A2 (new_n7587_),
	   .A1 (new_n7585_) );
   BUF_X4 g0857 (
	   .Z (new_n7587_),
	   .A (new_n7586_1_) );
   NOR2_X1 g0856 (
	   .ZN (new_n7586_1_),
	   .A2 (new_n7552_),
	   .A1 (new_n7200_) );
   NAND4_X1 g0855 (
	   .ZN (new_n7585_),
	   .A4 (new_n7584_),
	   .A3 (new_n7583_),
	   .A2 (new_n7582_),
	   .A1 (new_n7581_1_) );
   NAND3_X1 g0854 (
	   .ZN (new_n7584_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6804) );
   NAND3_X1 g0853 (
	   .ZN (new_n7583_),
	   .A3 (net_6772),
	   .A2 (_net_6824),
	   .A1 (new_n7570_) );
   NAND3_X1 g0852 (
	   .ZN (new_n7582_),
	   .A3 (_net_6823),
	   .A2 (net_6740),
	   .A1 (new_n7568_) );
   NAND2_X1 g0851 (
	   .ZN (new_n7581_1_),
	   .A2 (net_6708),
	   .A1 (new_n7566_) );
   NAND2_X1 g0850 (
	   .ZN (new_n7580_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n7579_) );
   NAND4_X1 g0849 (
	   .ZN (new_n7579_),
	   .A4 (new_n7578_),
	   .A3 (new_n7577_1_),
	   .A2 (new_n7576_),
	   .A1 (new_n7575_) );
   NAND3_X1 g0848 (
	   .ZN (new_n7578_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6806) );
   NAND3_X1 g0847 (
	   .ZN (new_n7577_1_),
	   .A3 (_net_6824),
	   .A2 (net_6774),
	   .A1 (new_n7570_) );
   NAND3_X1 g0846 (
	   .ZN (new_n7576_),
	   .A3 (net_6742),
	   .A2 (_net_6823),
	   .A1 (new_n7568_) );
   NAND2_X1 g0845 (
	   .ZN (new_n7575_),
	   .A2 (net_6710),
	   .A1 (new_n7566_) );
   NAND2_X1 g0844 (
	   .ZN (new_n7574_),
	   .A2 (new_n7573_),
	   .A1 (new_n7565_) );
   NAND4_X1 g0843 (
	   .ZN (new_n7573_),
	   .A4 (new_n7572_1_),
	   .A3 (new_n7571_),
	   .A2 (new_n7569_),
	   .A1 (new_n7567_1_) );
   NAND3_X1 g0842 (
	   .ZN (new_n7572_1_),
	   .A3 (_net_6824),
	   .A2 (_net_6823),
	   .A1 (net_6802) );
   NAND3_X1 g0841 (
	   .ZN (new_n7571_),
	   .A3 (_net_6824),
	   .A2 (net_6770),
	   .A1 (new_n7570_) );
   BUF_X4 g0840 (
	   .Z (new_n7570_),
	   .A (new_n7186_) );
   NAND3_X1 g0839 (
	   .ZN (new_n7569_),
	   .A3 (_net_6823),
	   .A2 (net_6738),
	   .A1 (new_n7568_) );
   BUF_X4 g0838 (
	   .Z (new_n7568_),
	   .A (new_n7187_) );
   NAND2_X1 g0837 (
	   .ZN (new_n7567_1_),
	   .A2 (net_6706),
	   .A1 (new_n7566_) );
   BUF_X4 g0836 (
	   .Z (new_n7566_),
	   .A (new_n7195_) );
   BUF_X4 g0835 (
	   .Z (new_n7565_),
	   .A (new_n7564_) );
   NOR3_X1 g0834 (
	   .ZN (new_n7564_),
	   .A3 (_net_6822),
	   .A2 (new_n7553_1_),
	   .A1 (new_n7200_) );
   AND4_X1 g0833 (
	   .ZN (new_n7563_1_),
	   .A4 (new_n7562_),
	   .A3 (new_n7561_),
	   .A2 (new_n7558_1_),
	   .A1 (new_n7557_) );
   NAND4_X1 g0832 (
	   .ZN (new_n7562_),
	   .A4 (new_n7194_1_),
	   .A3 (net_6754),
	   .A2 (_net_6822),
	   .A1 (new_n7560_) );
   NAND4_X1 g0831 (
	   .ZN (new_n7561_),
	   .A4 (new_n7191_),
	   .A3 (net_6786),
	   .A2 (_net_6822),
	   .A1 (new_n7560_) );
   BUF_X4 g0830 (
	   .Z (new_n7560_),
	   .A (new_n7559_) );
   NOR2_X2 g0829 (
	   .ZN (new_n7559_),
	   .A2 (new_n7553_1_),
	   .A1 (new_n7200_) );
   NAND3_X1 g0828 (
	   .ZN (new_n7558_1_),
	   .A3 (new_n7189_),
	   .A2 (net_6818),
	   .A1 (new_n7555_) );
   NAND3_X1 g0827 (
	   .ZN (new_n7557_),
	   .A3 (new_n7196_),
	   .A2 (net_6722),
	   .A1 (new_n7556_) );
   BUF_X4 g0826 (
	   .Z (new_n7556_),
	   .A (new_n7555_) );
   NOR3_X2 g0825 (
	   .ZN (new_n7555_),
	   .A3 (new_n7554_),
	   .A2 (new_n7553_1_),
	   .A1 (new_n7200_) );
   INV_X1 g0824 (
	   .ZN (new_n7554_),
	   .A (_net_6822) );
   NAND2_X1 g0823 (
	   .ZN (new_n7553_1_),
	   .A2 (new_n7201_),
	   .A1 (new_n7552_) );
   INV_X1 g0822 (
	   .ZN (new_n7552_),
	   .A (_net_6008) );
   MUX2_X1 g0821 (
	   .Z (n1010),
	   .S (new_n7504_),
	   .B (_net_7621),
	   .A (new_n7542_) );
   CLKBUF_X1 g0820 (
	   .Z (n1005),
	   .A (net_6391) );
   CLKBUF_X1 g0819 (
	   .Z (n1000),
	   .A (net_388) );
   NOR2_X1 g0818 (
	   .ZN (n995),
	   .A2 (x1006),
	   .A1 (new_n7547_) );
   AOI21_X1 g0817 (
	   .ZN (new_n7547_),
	   .B2 (net_7774),
	   .B1 (new_n7345_),
	   .A (_net_5856) );
   MUX2_X1 g0816 (
	   .Z (n990),
	   .S (new_n7545_),
	   .B (_net_7653),
	   .A (new_n7542_) );
   BUF_X8 g0815 (
	   .Z (new_n7545_),
	   .A (new_n7544_) );
   NAND2_X1 g0814 (
	   .ZN (new_n7544_),
	   .A2 (new_n7543_1_),
	   .A1 (new_n7026_) );
   NOR2_X1 g0813 (
	   .ZN (new_n7543_1_),
	   .A2 (new_n7027_1_),
	   .A1 (new_n7502_) );
   OAI21_X1 g0812 (
	   .ZN (new_n7542_),
	   .B2 (new_n7541_),
	   .B1 (new_n7020_),
	   .A (new_n7540_) );
   INV_X1 g0811 (
	   .ZN (new_n7541_),
	   .A (net_7541) );
   AOI22_X1 g0810 (
	   .ZN (new_n7540_),
	   .B2 (_net_291),
	   .B1 (net_373),
	   .A2 (_net_292),
	   .A1 (net_371) );
   MUX2_X1 g0809 (
	   .Z (n985),
	   .S (new_n7538_),
	   .B (_net_282),
	   .A (_net_7805) );
   BUF_X8 g0808 (
	   .Z (new_n7538_),
	   .A (new_n7537_) );
   NAND2_X2 g0807 (
	   .ZN (new_n7537_),
	   .A2 (new_n6820_),
	   .A1 (new_n7283_) );
   CLKBUF_X1 g0806 (
	   .Z (n981),
	   .A (net_6999) );
   CLKBUF_X1 g0805 (
	   .Z (n976),
	   .A (_net_7813) );
   OAI21_X1 g0804 (
	   .ZN (n971),
	   .B2 (new_n7258_),
	   .B1 (new_n7533_),
	   .A (new_n7532_) );
   INV_X1 g0803 (
	   .ZN (new_n7533_),
	   .A (_net_7296) );
   NAND2_X1 g0802 (
	   .ZN (new_n7532_),
	   .A2 (new_n7531_),
	   .A1 (new_n7252_1_) );
   OAI21_X1 g0801 (
	   .ZN (new_n7531_),
	   .B2 (new_n7530_1_),
	   .B1 (new_n6952_1_),
	   .A (new_n7529_) );
   INV_X1 g0800 (
	   .ZN (new_n7530_1_),
	   .A (net_7248) );
   AOI22_X1 g0799 (
	   .ZN (new_n7529_),
	   .B2 (net_342),
	   .B1 (_net_269),
	   .A2 (net_340),
	   .A1 (_net_270) );
   OAI221_X1 g0798 (
	   .ZN (n966),
	   .C2 (new_n7303_),
	   .C1 (new_n7527_1_),
	   .B2 (new_n7306_),
	   .B1 (new_n7526_),
	   .A (new_n7525_) );
   INV_X1 g0797 (
	   .ZN (new_n7527_1_),
	   .A (_net_7476) );
   INV_X1 g0796 (
	   .ZN (new_n7526_),
	   .A (_net_7508) );
   AOI22_X1 g0795 (
	   .ZN (new_n7525_),
	   .B2 (_net_7412),
	   .B1 (new_n7298_),
	   .A2 (_net_7444),
	   .A1 (new_n7296_) );
   MUX2_X1 g0794 (
	   .Z (n961),
	   .S (new_n7504_),
	   .B (_net_7629),
	   .A (new_n7523_) );
   OAI21_X1 g0793 (
	   .ZN (new_n7523_),
	   .B2 (new_n7522_1_),
	   .B1 (new_n7020_),
	   .A (new_n7521_) );
   INV_X1 g0792 (
	   .ZN (new_n7522_1_),
	   .A (net_7549) );
   AOI22_X1 g0791 (
	   .ZN (new_n7521_),
	   .B2 (_net_292),
	   .B1 (net_379),
	   .A2 (_net_291),
	   .A1 (net_381) );
   CLKBUF_X1 g0790 (
	   .Z (n956),
	   .A (_net_7823) );
   CLKBUF_X1 g0789 (
	   .Z (n953),
	   .A (net_6989) );
   CLKBUF_X1 g0788 (
	   .Z (n948),
	   .A (x1467) );
   AOI21_X1 g0787 (
	   .ZN (n944),
	   .B2 (new_n7516_),
	   .B1 (new_n7515_),
	   .A (x868) );
   INV_X1 g0786 (
	   .ZN (new_n7516_),
	   .A (_net_5851) );
   NAND3_X1 g0785 (
	   .ZN (new_n7515_),
	   .A3 (_net_284),
	   .A2 (net_7779),
	   .A1 (n3827) );
   AOI21_X1 g0784 (
	   .ZN (n3827),
	   .B2 (new_n7513_1_),
	   .B1 (new_n7512_),
	   .A (new_n7508_) );
   AOI21_X1 g0783 (
	   .ZN (new_n7513_1_),
	   .B2 (new_n7511_),
	   .B1 (new_n7510_),
	   .A (_net_226) );
   OAI21_X1 g0782 (
	   .ZN (new_n7512_),
	   .B2 (new_n7511_),
	   .B1 (new_n7510_),
	   .A (new_n7509_1_) );
   INV_X1 g0781 (
	   .ZN (new_n7511_),
	   .A (_net_229) );
   NOR2_X1 g0780 (
	   .ZN (new_n7510_),
	   .A2 (_net_228),
	   .A1 (_net_282) );
   INV_X1 g0779 (
	   .ZN (new_n7509_1_),
	   .A (_net_283) );
   INV_X1 g0778 (
	   .ZN (new_n7508_),
	   .A (_net_278) );
   CLKBUF_X1 g0777 (
	   .Z (n940),
	   .A (net_6979) );
   CLKBUF_X1 g0776 (
	   .Z (n935),
	   .A (net_7799) );
   MUX2_X1 g0775 (
	   .Z (n930),
	   .S (new_n7504_),
	   .B (_net_7632),
	   .A (new_n7501_1_) );
   BUF_X8 g0774 (
	   .Z (new_n7504_),
	   .A (new_n7503_) );
   NAND3_X1 g0773 (
	   .ZN (new_n7503_),
	   .A3 (_net_7685),
	   .A2 (new_n7502_),
	   .A1 (new_n7026_) );
   INV_X1 g0772 (
	   .ZN (new_n7502_),
	   .A (_net_7684) );
   OAI21_X1 g0771 (
	   .ZN (new_n7501_1_),
	   .B2 (new_n7500_),
	   .B1 (new_n7020_),
	   .A (new_n7499_) );
   INV_X1 g0770 (
	   .ZN (new_n7500_),
	   .A (net_370) );
   AOI22_X1 g0769 (
	   .ZN (new_n7499_),
	   .B2 (net_384),
	   .B1 (_net_291),
	   .A2 (_net_292),
	   .A1 (net_382) );
   OAI21_X1 g0768 (
	   .ZN (n925),
	   .B2 (new_n7111_1_),
	   .B1 (new_n7497_),
	   .A (new_n7496_1_) );
   INV_X1 g0767 (
	   .ZN (new_n7497_),
	   .A (_net_7354) );
   NAND2_X1 g0766 (
	   .ZN (new_n7496_1_),
	   .A2 (new_n7495_),
	   .A1 (new_n7101_) );
   OAI221_X1 g0765 (
	   .ZN (new_n7495_),
	   .C2 (new_n7105_),
	   .C1 (new_n7494_),
	   .B2 (new_n7106_),
	   .B1 (new_n7493_),
	   .A (new_n7492_1_) );
   INV_X1 g0764 (
	   .ZN (new_n7494_),
	   .A (net_336) );
   INV_X1 g0763 (
	   .ZN (new_n7493_),
	   .A (net_334) );
   NAND2_X1 g0762 (
	   .ZN (new_n7492_1_),
	   .A2 (net_7242),
	   .A1 (new_n7102_1_) );
   CLKBUF_X1 g0761 (
	   .Z (n920),
	   .A (_net_6160) );
   CLKBUF_X1 g0760 (
	   .Z (n916),
	   .A (net_6746) );
   CLKBUF_X1 g0759 (
	   .Z (n911),
	   .A (_net_7806) );
   CLKBUF_X1 g0758 (
	   .Z (n907),
	   .A (_net_7800) );
   OAI21_X1 g0757 (
	   .ZN (n903),
	   .B2 (new_n7279_),
	   .B1 (new_n7486_),
	   .A (new_n7485_) );
   INV_X1 g0756 (
	   .ZN (new_n7486_),
	   .A (_net_7439) );
   NAND2_X1 g0755 (
	   .ZN (new_n7485_),
	   .A2 (new_n7484_),
	   .A1 (new_n7272_) );
   OAI221_X1 g0754 (
	   .ZN (new_n7484_),
	   .C2 (new_n7275_1_),
	   .C1 (new_n6902_1_),
	   .B2 (new_n6901_),
	   .B1 (new_n7483_),
	   .A (new_n7482_1_) );
   INV_X1 g0753 (
	   .ZN (new_n7483_),
	   .A (net_352) );
   NAND2_X1 g0752 (
	   .ZN (new_n7482_1_),
	   .A2 (net_7391),
	   .A1 (new_n6898_) );
   CLKBUF_X1 g0751 (
	   .Z (n899),
	   .A (net_6739) );
   CLKBUF_X1 g0750 (
	   .Z (n894),
	   .A (net_6382) );
   CLKBUF_X1 g0749 (
	   .Z (n890),
	   .A (net_6616) );
   MUX2_X1 g0748 (
	   .Z (n885),
	   .S (new_n7437_1_),
	   .B (_net_6008),
	   .A (_net_7811) );
   CLKBUF_X1 g0747 (
	   .Z (n880),
	   .A (_net_7816) );
   NOR2_X1 g0746 (
	   .ZN (n875),
	   .A2 (new_n7334_),
	   .A1 (new_n6952_1_) );
   CLKBUF_X1 g0745 (
	   .Z (n870),
	   .A (_net_7818) );
   CLKBUF_X1 g0744 (
	   .Z (n867),
	   .A (net_6711) );
   NAND2_X1 g0743 (
	   .ZN (n862),
	   .A2 (new_n7472_),
	   .A1 (new_n7471_) );
   NAND2_X1 g0742 (
	   .ZN (new_n7472_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n7011_) );
   AOI22_X1 g0741 (
	   .ZN (new_n7471_),
	   .B2 (new_n6985_),
	   .B1 (_net_6086),
	   .A2 (new_n6980_),
	   .A1 (new_n6992_) );
   CLKBUF_X1 g0740 (
	   .Z (n857),
	   .A (_net_7794) );
   CLKBUF_X1 g0739 (
	   .Z (n854),
	   .A (net_7390) );
   OAI221_X1 g0738 (
	   .ZN (n849),
	   .C2 (new_n6920_),
	   .C1 (new_n7467_),
	   .B2 (new_n6917_),
	   .B1 (new_n7466_),
	   .A (new_n7465_) );
   INV_X1 g0737 (
	   .ZN (new_n7467_),
	   .A (_net_7361) );
   INV_X1 g0736 (
	   .ZN (new_n7466_),
	   .A (_net_7297) );
   AOI22_X1 g0735 (
	   .ZN (new_n7465_),
	   .B2 (_net_7265),
	   .B1 (new_n6913_),
	   .A2 (_net_7329),
	   .A1 (new_n6911_) );
   CLKBUF_X1 g0734 (
	   .Z (n844),
	   .A (net_6381) );
   CLKBUF_X1 g0733 (
	   .Z (n839),
	   .A (_net_7818) );
   NAND2_X1 g0732 (
	   .ZN (n834),
	   .A2 (new_n7461_),
	   .A1 (new_n7459_1_) );
   AOI22_X1 g0731 (
	   .ZN (new_n7461_),
	   .B2 (net_7524),
	   .B1 (new_n7460_),
	   .A2 (new_n7301_),
	   .A1 (net_7492) );
   INV_X2 g0730 (
	   .ZN (new_n7460_),
	   .A (new_n7305_) );
   AOI22_X1 g0729 (
	   .ZN (new_n7459_1_),
	   .B2 (_net_7428),
	   .B1 (new_n7298_),
	   .A2 (net_7460),
	   .A1 (new_n7296_) );
   CLKBUF_X1 g0728 (
	   .Z (n830),
	   .A (net_7396) );
   MUX2_X1 g0727 (
	   .Z (n825),
	   .S (_net_154),
	   .B (net_316),
	   .A (_net_120) );
   MUX2_X1 g0726 (
	   .Z (n820),
	   .S (_net_154),
	   .B (net_317),
	   .A (_net_121) );
   CLKBUF_X1 g0725 (
	   .Z (n815),
	   .A (_net_6084) );
   CLKBUF_X1 g0724 (
	   .Z (n811),
	   .A (net_6399) );
   NOR3_X1 g0723 (
	   .ZN (n806),
	   .A3 (new_n7452_),
	   .A2 (new_n7451_),
	   .A1 (new_n7449_) );
   AOI21_X1 g0722 (
	   .ZN (new_n7452_),
	   .B2 (_net_7784),
	   .B1 (_net_7785),
	   .A (_net_7786) );
   INV_X1 g0721 (
	   .ZN (new_n7451_),
	   .A (new_n7450_1_) );
   NAND3_X1 g0720 (
	   .ZN (new_n7450_1_),
	   .A3 (_net_7784),
	   .A2 (_net_7785),
	   .A1 (_net_7786) );
   INV_X1 g0719 (
	   .ZN (new_n7449_),
	   .A (new_n7448_) );
   NOR2_X1 g0718 (
	   .ZN (new_n7448_),
	   .A2 (_net_113),
	   .A1 (new_n7447_) );
   NOR2_X1 g0717 (
	   .ZN (new_n7447_),
	   .A2 (new_n7446_1_),
	   .A1 (new_n7444_) );
   NAND2_X1 g0716 (
	   .ZN (new_n7446_1_),
	   .A2 (_net_7784),
	   .A1 (new_n7445_) );
   INV_X1 g0715 (
	   .ZN (new_n7445_),
	   .A (_net_7785) );
   NAND4_X1 g0714 (
	   .ZN (new_n7444_),
	   .A4 (_net_7788),
	   .A3 (_net_7789),
	   .A2 (new_n7443_),
	   .A1 (new_n7442_1_) );
   INV_X1 g0713 (
	   .ZN (new_n7443_),
	   .A (_net_7787) );
   INV_X1 g0712 (
	   .ZN (new_n7442_1_),
	   .A (_net_7786) );
   CLKBUF_X1 g0711 (
	   .Z (n802),
	   .A (net_7133) );
   CLKBUF_X1 g0710 (
	   .Z (n798),
	   .A (net_7134) );
   AND2_X1 g0709 (
	   .ZN (n793),
	   .A2 (net_377),
	   .A1 (new_n7262_) );
   MUX2_X1 g0708 (
	   .Z (n788),
	   .S (new_n7437_1_),
	   .B (_net_6012),
	   .A (_net_7815) );
   BUF_X8 g0707 (
	   .Z (new_n7437_1_),
	   .A (new_n7436_) );
   BUF_X8 g0706 (
	   .Z (new_n7436_),
	   .A (new_n7435_) );
   NAND2_X1 g0705 (
	   .ZN (new_n7435_),
	   .A2 (new_n7364_),
	   .A1 (new_n7283_) );
   CLKBUF_X1 g0704 (
	   .Z (n783),
	   .A (net_7802) );
   CLKBUF_X1 g0703 (
	   .Z (n779),
	   .A (net_6385) );
   CLKBUF_X1 g0702 (
	   .Z (n774),
	   .A (x806) );
   AOI21_X1 g0701 (
	   .ZN (n770),
	   .B2 (new_n7430_),
	   .B1 (new_n7429_),
	   .A (new_n7428_) );
   INV_X1 g0700 (
	   .ZN (new_n7430_),
	   .A (_net_6026) );
   INV_X1 g0699 (
	   .ZN (new_n7429_),
	   .A (_net_7732) );
   BUF_X4 g0698 (
	   .Z (new_n7428_),
	   .A (new_n7427_1_) );
   INV_X1 g0697 (
	   .ZN (new_n7427_1_),
	   .A (n1792) );
   NAND2_X1 g0696 (
	   .ZN (n1792),
	   .A2 (n4304),
	   .A1 (new_n7422_1_) );
   NOR2_X2 g0695 (
	   .ZN (n4304),
	   .A2 (new_n7177_1_),
	   .A1 (new_n7424_) );
   NAND3_X1 g0694 (
	   .ZN (new_n7424_),
	   .A3 (_net_7687),
	   .A2 (new_n7423_),
	   .A1 (new_n7178_) );
   INV_X1 g0693 (
	   .ZN (new_n7423_),
	   .A (_net_7688) );
   AND3_X2 g0692 (
	   .ZN (new_n7422_1_),
	   .A3 (new_n7394_),
	   .A2 (new_n7356_),
	   .A1 (new_n7392_) );
   AND3_X1 g0691 (
	   .ZN (n765),
	   .A3 (new_n7364_),
	   .A2 (_net_7793),
	   .A1 (new_n6822_1_) );
   CLKBUF_X1 g0690 (
	   .Z (n761),
	   .A (net_6468) );
   NAND2_X1 g0689 (
	   .ZN (n756),
	   .A2 (new_n7418_),
	   .A1 (new_n7414_) );
   NAND2_X1 g0688 (
	   .ZN (new_n7418_),
	   .A2 (new_n7070_),
	   .A1 (new_n7417_1_) );
   NAND2_X1 g0687 (
	   .ZN (new_n7417_1_),
	   .A2 (new_n7416_),
	   .A1 (new_n7415_) );
   AOI22_X1 g0686 (
	   .ZN (new_n7416_),
	   .B2 (net_6965),
	   .B1 (new_n7052_),
	   .A2 (net_6997),
	   .A1 (new_n7050_) );
   AOI22_X1 g0685 (
	   .ZN (new_n7415_),
	   .B2 (net_7061),
	   .B1 (new_n7046_),
	   .A2 (new_n7044_),
	   .A1 (net_7029) );
   AOI22_X1 g0684 (
	   .ZN (new_n7414_),
	   .B2 (new_n7092_),
	   .B1 (_net_6147),
	   .A2 (new_n7089_1_),
	   .A1 (new_n7413_1_) );
   NAND2_X1 g0683 (
	   .ZN (new_n7413_1_),
	   .A2 (new_n7412_),
	   .A1 (new_n7411_) );
   AOI22_X1 g0682 (
	   .ZN (new_n7412_),
	   .B2 (net_6967),
	   .B1 (new_n7052_),
	   .A2 (net_6999),
	   .A1 (new_n7050_) );
   AOI22_X1 g0681 (
	   .ZN (new_n7411_),
	   .B2 (net_7063),
	   .B1 (new_n7046_),
	   .A2 (new_n7044_),
	   .A1 (net_7031) );
   CLKBUF_X1 g0680 (
	   .Z (n751),
	   .A (_net_5976) );
   NAND2_X1 g0679 (
	   .ZN (n746),
	   .A2 (new_n7408_1_),
	   .A1 (new_n7407_) );
   AOI22_X1 g0678 (
	   .ZN (new_n7408_1_),
	   .B2 (_net_7557),
	   .B1 (new_n6755_),
	   .A2 (_net_7621),
	   .A1 (new_n6746_1_) );
   AOI22_X1 g0677 (
	   .ZN (new_n7407_),
	   .B2 (_net_7589),
	   .B1 (new_n7350_),
	   .A2 (new_n6749_1_),
	   .A1 (_net_7653) );
   CLKBUF_X1 g0676 (
	   .Z (n741),
	   .A (net_147) );
   NAND2_X1 g0675 (
	   .ZN (n736),
	   .A2 (new_n7404_1_),
	   .A1 (new_n7403_) );
   INV_X1 g0674 (
	   .ZN (new_n7404_1_),
	   .A (_net_6037) );
   NAND2_X1 g0673 (
	   .ZN (new_n7403_),
	   .A2 (_net_5976),
	   .A1 (new_n7056_) );
   NAND3_X1 g0672 (
	   .ZN (n732),
	   .A3 (new_n7401_),
	   .A2 (new_n7398_),
	   .A1 (new_n7368_1_) );
   NAND4_X1 g0671 (
	   .ZN (new_n7401_),
	   .A4 (_net_7701),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n7400_1_) );
   BUF_X4 g0670 (
	   .Z (new_n7400_1_),
	   .A (new_n7399_) );
   AND2_X2 g0669 (
	   .ZN (new_n7399_),
	   .A2 (new_n7360_),
	   .A1 (new_n7357_) );
   NOR3_X1 g0668 (
	   .ZN (new_n7398_),
	   .A3 (new_n7397_),
	   .A2 (new_n7379_),
	   .A1 (new_n7372_1_) );
   NAND3_X1 g0667 (
	   .ZN (new_n7397_),
	   .A3 (new_n7396_),
	   .A2 (new_n7390_),
	   .A1 (new_n7384_) );
   NAND4_X1 g0666 (
	   .ZN (new_n7396_),
	   .A4 (net_166),
	   .A3 (x1231),
	   .A2 (new_n7395_1_),
	   .A1 (new_n7393_) );
   BUF_X4 g0665 (
	   .Z (new_n7395_1_),
	   .A (new_n7394_) );
   NOR2_X2 g0664 (
	   .ZN (new_n7394_),
	   .A2 (x1215),
	   .A1 (x1322) );
   BUF_X4 g0663 (
	   .Z (new_n7393_),
	   .A (new_n7392_) );
   BUF_X4 g0662 (
	   .Z (new_n7392_),
	   .A (new_n7391_1_) );
   AND2_X1 g0661 (
	   .ZN (new_n7391_1_),
	   .A2 (x1286),
	   .A1 (x1261) );
   NAND3_X1 g0660 (
	   .ZN (new_n7390_),
	   .A3 (net_203),
	   .A2 (new_n7389_),
	   .A1 (new_n7387_) );
   BUF_X4 g0659 (
	   .Z (new_n7389_),
	   .A (new_n7388_) );
   NOR2_X2 g0658 (
	   .ZN (new_n7388_),
	   .A2 (x1215),
	   .A1 (new_n7282_) );
   BUF_X4 g0657 (
	   .Z (new_n7387_),
	   .A (new_n7386_1_) );
   BUF_X4 g0656 (
	   .Z (new_n7386_1_),
	   .A (new_n7385_) );
   AND3_X1 g0655 (
	   .ZN (new_n7385_),
	   .A3 (x1231),
	   .A2 (x1286),
	   .A1 (x1261) );
   NAND3_X1 g0654 (
	   .ZN (new_n7384_),
	   .A3 (net_240),
	   .A2 (new_n7383_),
	   .A1 (new_n7381_1_) );
   BUF_X4 g0653 (
	   .Z (new_n7383_),
	   .A (new_n7382_) );
   NOR2_X2 g0652 (
	   .ZN (new_n7382_),
	   .A2 (x1231),
	   .A1 (new_n7358_) );
   BUF_X4 g0651 (
	   .Z (new_n7381_1_),
	   .A (new_n7380_) );
   NOR3_X2 g0650 (
	   .ZN (new_n7380_),
	   .A3 (x1286),
	   .A2 (x1261),
	   .A1 (x1322) );
   OAI22_X1 g0649 (
	   .ZN (new_n7379_),
	   .B2 (new_n7378_),
	   .B1 (new_n7376_1_),
	   .A2 (new_n7375_),
	   .A1 (new_n7374_) );
   BUF_X4 g0648 (
	   .Z (new_n7378_),
	   .A (new_n7377_) );
   OAI211_X1 g0647 (
	   .ZN (new_n7377_),
	   .C2 (x1215),
	   .C1 (new_n7356_),
	   .B (x1286),
	   .A (x1261) );
   INV_X1 g0646 (
	   .ZN (new_n7376_1_),
	   .A (_net_7730) );
   INV_X1 g0645 (
	   .ZN (new_n7375_),
	   .A (_net_124) );
   OAI211_X2 g0644 (
	   .ZN (new_n7374_),
	   .C2 (x1215),
	   .C1 (new_n7373_),
	   .B (new_n7354_1_),
	   .A (x1261) );
   NAND3_X1 g0643 (
	   .ZN (new_n7373_),
	   .A3 (x1231),
	   .A2 (x1286),
	   .A1 (x1261) );
   AND4_X1 g0642 (
	   .ZN (new_n7372_1_),
	   .A4 (new_n7371_),
	   .A3 (new_n7370_),
	   .A2 (new_n7369_),
	   .A1 (_net_6041) );
   NOR3_X2 g0641 (
	   .ZN (new_n7371_),
	   .A3 (x1261),
	   .A2 (x1322),
	   .A1 (new_n6819_) );
   BUF_X4 g0640 (
	   .Z (new_n7370_),
	   .A (new_n7360_) );
   BUF_X4 g0639 (
	   .Z (new_n7369_),
	   .A (new_n7357_) );
   NOR2_X1 g0638 (
	   .ZN (new_n7368_1_),
	   .A2 (new_n7367_),
	   .A1 (new_n7363_1_) );
   NOR2_X1 g0637 (
	   .ZN (new_n7367_),
	   .A2 (new_n6993_),
	   .A1 (new_n7366_) );
   BUF_X4 g0636 (
	   .Z (new_n7366_),
	   .A (new_n7365_) );
   NAND4_X1 g0635 (
	   .ZN (new_n7365_),
	   .A4 (new_n7364_),
	   .A3 (new_n7359_1_),
	   .A2 (x1322),
	   .A1 (new_n7357_) );
   NOR2_X2 g0634 (
	   .ZN (new_n7364_),
	   .A2 (x1286),
	   .A1 (x1261) );
   NOR2_X1 g0633 (
	   .ZN (new_n7363_1_),
	   .A2 (new_n6902_1_),
	   .A1 (new_n7362_) );
   BUF_X4 g0632 (
	   .Z (new_n7362_),
	   .A (new_n7361_) );
   NAND4_X1 g0631 (
	   .ZN (new_n7361_),
	   .A4 (new_n7360_),
	   .A3 (x1286),
	   .A2 (x1322),
	   .A1 (new_n7357_) );
   BUF_X4 g0630 (
	   .Z (new_n7360_),
	   .A (new_n7359_1_) );
   NAND4_X1 g0629 (
	   .ZN (new_n7359_1_),
	   .A4 (x1231),
	   .A3 (x1286),
	   .A2 (x1261),
	   .A1 (new_n7358_) );
   INV_X1 g0628 (
	   .ZN (new_n7358_),
	   .A (x1215) );
   NAND4_X1 g0627 (
	   .ZN (new_n7357_),
	   .A4 (new_n7356_),
	   .A3 (new_n7355_),
	   .A2 (x1215),
	   .A1 (new_n7354_1_) );
   INV_X1 g0626 (
	   .ZN (new_n7356_),
	   .A (x1231) );
   INV_X1 g0625 (
	   .ZN (new_n7355_),
	   .A (x1261) );
   NOR2_X2 g0624 (
	   .ZN (new_n7354_1_),
	   .A2 (x1286),
	   .A1 (x1322) );
   NAND2_X1 g0623 (
	   .ZN (n727),
	   .A2 (new_n7352_),
	   .A1 (new_n7351_) );
   AOI22_X1 g0622 (
	   .ZN (new_n7352_),
	   .B2 (_net_7558),
	   .B1 (new_n6755_),
	   .A2 (_net_7622),
	   .A1 (new_n6746_1_) );
   AOI22_X1 g0621 (
	   .ZN (new_n7351_),
	   .B2 (_net_7590),
	   .B1 (new_n7350_),
	   .A2 (new_n6749_1_),
	   .A1 (_net_7654) );
   BUF_X4 g0620 (
	   .Z (new_n7350_),
	   .A (new_n6742_) );
   CLKBUF_X1 g0619 (
	   .Z (n722),
	   .A (net_6396) );
   AND2_X1 g0618 (
	   .ZN (n718),
	   .A2 (net_375),
	   .A1 (new_n7262_) );
   AND2_X1 g0617 (
	   .ZN (n713),
	   .A2 (new_n7346_),
	   .A1 (new_n7345_) );
   INV_X1 g0616 (
	   .ZN (new_n7346_),
	   .A (x1006) );
   AOI211_X1 g0615 (
	   .ZN (new_n7345_),
	   .C2 (new_n7344_1_),
	   .C1 (new_n7343_),
	   .B (new_n7208_),
	   .A (new_n7339_) );
   AOI21_X1 g0614 (
	   .ZN (new_n7344_1_),
	   .B2 (new_n7342_),
	   .B1 (new_n7341_),
	   .A (_net_5968) );
   OAI21_X1 g0613 (
	   .ZN (new_n7343_),
	   .B2 (new_n7342_),
	   .B1 (new_n7341_),
	   .A (new_n7340_1_) );
   INV_X1 g0612 (
	   .ZN (new_n7342_),
	   .A (_net_5970) );
   NOR2_X1 g0611 (
	   .ZN (new_n7341_),
	   .A2 (_net_6010),
	   .A1 (_net_5969) );
   INV_X1 g0610 (
	   .ZN (new_n7340_1_),
	   .A (_net_6011) );
   INV_X1 g0609 (
	   .ZN (new_n7339_),
	   .A (_net_6012) );
   OAI21_X1 g0608 (
	   .ZN (n708),
	   .B2 (new_n7258_),
	   .B1 (new_n7337_),
	   .A (new_n7336_) );
   INV_X1 g0607 (
	   .ZN (new_n7337_),
	   .A (_net_7300) );
   NAND2_X1 g0606 (
	   .ZN (new_n7336_),
	   .A2 (new_n7335_1_),
	   .A1 (new_n7252_1_) );
   OAI22_X1 g0605 (
	   .ZN (new_n7335_1_),
	   .B2 (new_n7334_),
	   .B1 (new_n7106_),
	   .A2 (new_n7333_),
	   .A1 (new_n6951_) );
   INV_X1 g0604 (
	   .ZN (new_n7334_),
	   .A (net_344) );
   INV_X1 g0603 (
	   .ZN (new_n7333_),
	   .A (net_332) );
   CLKBUF_X1 g0602 (
	   .Z (n703),
	   .A (_net_6127) );
   AND2_X1 g0601 (
	   .ZN (n698),
	   .A2 (net_383),
	   .A1 (new_n7262_) );
   AOI21_X1 g0600 (
	   .ZN (n693),
	   .B2 (new_n7326_1_),
	   .B1 (new_n7329_),
	   .A (new_n7328_) );
   INV_X1 g0599 (
	   .ZN (new_n7329_),
	   .A (_net_7271) );
   NOR2_X1 g0598 (
	   .ZN (new_n7328_),
	   .A2 (n1350),
	   .A1 (new_n7326_1_) );
   NOR2_X1 g0597 (
	   .ZN (n1350),
	   .A2 (new_n7107_1_),
	   .A1 (new_n6952_1_) );
   BUF_X4 g0596 (
	   .Z (new_n7326_1_),
	   .A (new_n7325_) );
   NAND2_X2 g0595 (
	   .ZN (new_n7325_),
	   .A2 (new_n6946_),
	   .A1 (new_n6945_) );
   OAI21_X1 g0594 (
	   .ZN (n688),
	   .B2 (new_n7225_),
	   .B1 (new_n7323_),
	   .A (new_n7322_) );
   INV_X1 g0593 (
	   .ZN (new_n7323_),
	   .A (_net_7330) );
   NAND2_X1 g0592 (
	   .ZN (new_n7322_),
	   .A2 (new_n7321_1_),
	   .A1 (new_n7222_) );
   OAI21_X1 g0591 (
	   .ZN (new_n7321_1_),
	   .B2 (new_n7320_),
	   .B1 (new_n6952_1_),
	   .A (new_n7319_) );
   INV_X1 g0590 (
	   .ZN (new_n7320_),
	   .A (net_330) );
   AOI22_X1 g0589 (
	   .ZN (new_n7319_),
	   .B2 (net_344),
	   .B1 (_net_269),
	   .A2 (net_342),
	   .A1 (_net_270) );
   CLKBUF_X1 g0588 (
	   .Z (n683),
	   .A (_net_7796) );
   CLKBUF_X1 g0587 (
	   .Z (n678),
	   .A (_net_7823) );
   AND2_X1 g0586 (
	   .ZN (n673),
	   .A2 (_net_6207),
	   .A1 (new_n7239_) );
   CLKBUF_X1 g0585 (
	   .Z (n669),
	   .A (net_6440) );
   CLKBUF_X1 g0584 (
	   .Z (n664),
	   .A (net_6383) );
   OAI221_X1 g0583 (
	   .ZN (n659),
	   .C2 (new_n7312_1_),
	   .C1 (new_n7311_),
	   .B2 (new_n6920_),
	   .B1 (new_n7310_),
	   .A (new_n7309_) );
   BUF_X4 g0582 (
	   .Z (new_n7312_1_),
	   .A (new_n6916_) );
   INV_X1 g0581 (
	   .ZN (new_n7311_),
	   .A (_net_7286) );
   INV_X1 g0580 (
	   .ZN (new_n7310_),
	   .A (_net_7350) );
   AOI22_X1 g0579 (
	   .ZN (new_n7309_),
	   .B2 (_net_7254),
	   .B1 (new_n6913_),
	   .A2 (_net_7318),
	   .A1 (new_n6911_) );
   INV_X1 g0578 (
	   .ZN (n654),
	   .A (new_n7206_) );
   OAI221_X1 g0577 (
	   .ZN (n649),
	   .C2 (new_n7306_),
	   .C1 (new_n7304_),
	   .B2 (new_n7303_),
	   .B1 (new_n7300_),
	   .A (new_n7299_) );
   BUF_X4 g0576 (
	   .Z (new_n7306_),
	   .A (new_n7305_) );
   NAND2_X1 g0575 (
	   .ZN (new_n7305_),
	   .A2 (_net_7530),
	   .A1 (net_7529) );
   INV_X1 g0574 (
	   .ZN (new_n7304_),
	   .A (_net_7516) );
   BUF_X4 g0573 (
	   .Z (new_n7303_),
	   .A (new_n7302_1_) );
   INV_X1 g0572 (
	   .ZN (new_n7302_1_),
	   .A (new_n7301_) );
   NOR2_X2 g0571 (
	   .ZN (new_n7301_),
	   .A2 (net_7529),
	   .A1 (new_n7294_) );
   INV_X1 g0570 (
	   .ZN (new_n7300_),
	   .A (_net_7484) );
   AOI22_X1 g0569 (
	   .ZN (new_n7299_),
	   .B2 (_net_7420),
	   .B1 (new_n7298_),
	   .A2 (_net_7452),
	   .A1 (new_n7296_) );
   BUF_X4 g0568 (
	   .Z (new_n7298_),
	   .A (new_n7297_1_) );
   NOR2_X1 g0567 (
	   .ZN (new_n7297_1_),
	   .A2 (_net_7530),
	   .A1 (net_7529) );
   BUF_X4 g0566 (
	   .Z (new_n7296_),
	   .A (new_n7295_) );
   AND2_X1 g0565 (
	   .ZN (new_n7295_),
	   .A2 (net_7529),
	   .A1 (new_n7294_) );
   INV_X1 g0564 (
	   .ZN (new_n7294_),
	   .A (_net_7530) );
   OAI221_X1 g0563 (
	   .ZN (n644),
	   .C2 (new_n7292_1_),
	   .C1 (new_n7075_),
	   .B2 (new_n7291_),
	   .B1 (new_n7058_1_),
	   .A (new_n7288_1_) );
   INV_X1 g0562 (
	   .ZN (new_n7292_1_),
	   .A (new_n7092_) );
   NAND2_X1 g0561 (
	   .ZN (new_n7291_),
	   .A2 (new_n7290_),
	   .A1 (new_n7289_) );
   NAND3_X1 g0560 (
	   .ZN (new_n7290_),
	   .A3 (_net_7092),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   OAI21_X1 g0559 (
	   .ZN (new_n7289_),
	   .B2 (new_n7072_1_),
	   .B1 (new_n7077_1_),
	   .A (new_n7075_) );
   OAI21_X1 g0558 (
	   .ZN (new_n7288_1_),
	   .B2 (new_n7044_),
	   .B1 (new_n7050_),
	   .A (new_n7287_) );
   NOR2_X1 g0557 (
	   .ZN (new_n7287_),
	   .A2 (new_n7057_),
	   .A1 (new_n7067_1_) );
   MUX2_X1 g0556 (
	   .Z (n639),
	   .S (new_n7285_),
	   .B (_net_7694),
	   .A (_net_7796) );
   BUF_X8 g0555 (
	   .Z (new_n7285_),
	   .A (new_n7284_1_) );
   NAND3_X2 g0554 (
	   .ZN (new_n7284_1_),
	   .A3 (new_n6819_),
	   .A2 (x1261),
	   .A1 (new_n7283_) );
   NOR2_X1 g0553 (
	   .ZN (new_n7283_),
	   .A2 (new_n6821_),
	   .A1 (new_n7282_) );
   INV_X1 g0552 (
	   .ZN (new_n7282_),
	   .A (x1322) );
   NOR2_X1 g0551 (
	   .ZN (n634),
	   .A2 (new_n7274_),
	   .A1 (new_n7035_) );
   OAI21_X1 g0550 (
	   .ZN (n629),
	   .B2 (new_n7279_),
	   .B1 (new_n7278_),
	   .A (new_n7277_) );
   BUF_X4 g0549 (
	   .Z (new_n7279_),
	   .A (new_n7271_) );
   INV_X1 g0548 (
	   .ZN (new_n7278_),
	   .A (_net_7441) );
   NAND2_X1 g0547 (
	   .ZN (new_n7277_),
	   .A2 (new_n7276_),
	   .A1 (new_n7272_) );
   OAI221_X1 g0546 (
	   .ZN (new_n7276_),
	   .C2 (new_n7275_1_),
	   .C1 (new_n6901_),
	   .B2 (new_n7274_),
	   .B1 (new_n6902_1_),
	   .A (new_n7273_) );
   INV_X1 g0545 (
	   .ZN (new_n7275_1_),
	   .A (net_354) );
   INV_X1 g0544 (
	   .ZN (new_n7274_),
	   .A (net_356) );
   NAND2_X1 g0543 (
	   .ZN (new_n7273_),
	   .A2 (net_7393),
	   .A1 (new_n6898_) );
   BUF_X4 g0542 (
	   .Z (new_n7272_),
	   .A (new_n7271_) );
   BUF_X4 g0541 (
	   .Z (new_n7271_),
	   .A (new_n7270_1_) );
   AND2_X1 g0540 (
	   .ZN (new_n7270_1_),
	   .A2 (new_n7269_),
	   .A1 (new_n6892_) );
   NOR2_X1 g0539 (
	   .ZN (new_n7269_),
	   .A2 (_net_7534),
	   .A1 (new_n7268_) );
   INV_X1 g0538 (
	   .ZN (new_n7268_),
	   .A (_net_7533) );
   CLKBUF_X1 g0537 (
	   .Z (n625),
	   .A (net_7246) );
   NAND2_X1 g0536 (
	   .ZN (n620),
	   .A2 (new_n7265_1_),
	   .A1 (new_n7264_) );
   INV_X1 g0535 (
	   .ZN (new_n7265_1_),
	   .A (_net_6004) );
   NAND2_X1 g0534 (
	   .ZN (new_n7264_),
	   .A2 (_net_5964),
	   .A1 (new_n6982_1_) );
   AND2_X1 g0533 (
	   .ZN (n615),
	   .A2 (net_374),
	   .A1 (new_n7262_) );
   BUF_X4 g0532 (
	   .Z (new_n7262_),
	   .A (new_n7018_1_) );
   CLKBUF_X1 g0531 (
	   .Z (n610),
	   .A (_net_7800) );
   AND2_X1 g0530 (
	   .ZN (n605),
	   .A2 (_net_6209),
	   .A1 (new_n7239_) );
   OAI21_X1 g0529 (
	   .ZN (n600),
	   .B2 (new_n7258_),
	   .B1 (new_n7257_),
	   .A (new_n7256_1_) );
   BUF_X4 g0528 (
	   .Z (new_n7258_),
	   .A (new_n7251_) );
   INV_X1 g0527 (
	   .ZN (new_n7257_),
	   .A (_net_7285) );
   NAND2_X1 g0526 (
	   .ZN (new_n7256_1_),
	   .A2 (new_n7255_),
	   .A1 (new_n7252_1_) );
   OAI21_X1 g0525 (
	   .ZN (new_n7255_),
	   .B2 (new_n7254_),
	   .B1 (new_n6952_1_),
	   .A (new_n7253_) );
   INV_X1 g0524 (
	   .ZN (new_n7254_),
	   .A (net_7237) );
   AOI22_X1 g0523 (
	   .ZN (new_n7253_),
	   .B2 (_net_269),
	   .B1 (net_331),
	   .A2 (_net_270),
	   .A1 (net_329) );
   BUF_X4 g0522 (
	   .Z (new_n7252_1_),
	   .A (new_n7251_) );
   BUF_X4 g0521 (
	   .Z (new_n7251_),
	   .A (new_n7250_) );
   AND2_X1 g0520 (
	   .ZN (new_n7250_),
	   .A2 (new_n7249_1_),
	   .A1 (new_n6945_) );
   NOR2_X1 g0519 (
	   .ZN (new_n7249_1_),
	   .A2 (_net_7383),
	   .A1 (new_n7248_) );
   INV_X1 g0518 (
	   .ZN (new_n7248_),
	   .A (_net_7382) );
   AND2_X1 g0517 (
	   .ZN (n595),
	   .A2 (net_361),
	   .A1 (new_n6898_) );
   CLKBUF_X1 g0516 (
	   .Z (n590),
	   .A (net_6400) );
   CLKBUF_X1 g0515 (
	   .Z (n585),
	   .A (_net_6177) );
   CLKBUF_X1 g0514 (
	   .Z (n580),
	   .A (x1587) );
   AND2_X1 g0513 (
	   .ZN (n576),
	   .A2 (net_342),
	   .A1 (new_n7102_1_) );
   CLKBUF_X1 g0512 (
	   .Z (n571),
	   .A (net_152) );
   CLKBUF_X1 g0511 (
	   .Z (n566),
	   .A (_net_7808) );
   AND2_X1 g0510 (
	   .ZN (n561),
	   .A2 (_net_6293),
	   .A1 (new_n7239_) );
   BUF_X2 g0509 (
	   .Z (new_n7239_),
	   .A (new_n7235_1_) );
   CLKBUF_X1 g0508 (
	   .Z (n556),
	   .A (_net_7794) );
   AOI21_X1 g0507 (
	   .ZN (n553),
	   .B2 (new_n7236_),
	   .B1 (new_n7234_),
	   .A (new_n7232_) );
   NOR3_X1 g0506 (
	   .ZN (new_n7236_),
	   .A3 (net_6058),
	   .A2 (net_6056),
	   .A1 (new_n7235_1_) );
   INV_X2 g0505 (
	   .ZN (new_n7235_1_),
	   .A (_net_392) );
   NOR3_X1 g0504 (
	   .ZN (new_n7234_),
	   .A3 (net_6060),
	   .A2 (_net_6062),
	   .A1 (new_n7233_) );
   OR4_X1 g0503 (
	   .ZN (new_n7233_),
	   .A4 (net_6061),
	   .A3 (net_6057),
	   .A2 (_net_6063),
	   .A1 (net_6059) );
   NOR2_X1 g0502 (
	   .ZN (new_n7232_),
	   .A2 (_net_392),
	   .A1 (_net_6199) );
   INV_X1 g0501 (
	   .ZN (n548),
	   .A (new_n7230_1_) );
   NAND2_X1 g0500 (
	   .ZN (new_n7230_1_),
	   .A2 (new_n7229_),
	   .A1 (new_n7227_) );
   NAND2_X1 g0499 (
	   .ZN (new_n7229_),
	   .A2 (_net_6688),
	   .A1 (new_n7228_) );
   INV_X1 g0498 (
	   .ZN (new_n7228_),
	   .A (net_6691) );
   NAND2_X1 g0497 (
	   .ZN (new_n7227_),
	   .A2 (net_6691),
	   .A1 (new_n7004_) );
   OAI21_X1 g0496 (
	   .ZN (n543),
	   .B2 (new_n7225_),
	   .B1 (new_n7224_),
	   .A (new_n7223_) );
   BUF_X4 g0495 (
	   .Z (new_n7225_),
	   .A (new_n7221_1_) );
   INV_X1 g0494 (
	   .ZN (new_n7224_),
	   .A (_net_7316) );
   NAND2_X1 g0493 (
	   .ZN (new_n7223_),
	   .A2 (new_n6954_),
	   .A1 (new_n7222_) );
   BUF_X4 g0492 (
	   .Z (new_n7222_),
	   .A (new_n7221_1_) );
   BUF_X4 g0491 (
	   .Z (new_n7221_1_),
	   .A (new_n7220_) );
   AND2_X1 g0490 (
	   .ZN (new_n7220_),
	   .A2 (new_n7219_),
	   .A1 (new_n6945_) );
   NOR2_X1 g0489 (
	   .ZN (new_n7219_),
	   .A2 (_net_7382),
	   .A1 (new_n7218_) );
   INV_X1 g0488 (
	   .ZN (new_n7218_),
	   .A (_net_7383) );
   MUX2_X1 g0487 (
	   .Z (n538),
	   .S (new_n7029_),
	   .B (_net_7603),
	   .A (new_n7216_1_) );
   OAI21_X1 g0486 (
	   .ZN (new_n7216_1_),
	   .B2 (new_n7215_),
	   .B1 (new_n7214_),
	   .A (new_n7213_) );
   INV_X1 g0485 (
	   .ZN (new_n7215_),
	   .A (_net_292) );
   INV_X1 g0484 (
	   .ZN (new_n7214_),
	   .A (net_385) );
   NAND2_X1 g0483 (
	   .ZN (new_n7213_),
	   .A2 (net_373),
	   .A1 (new_n7018_1_) );
   OAI21_X1 g0482 (
	   .ZN (n533),
	   .B2 (new_n7211_),
	   .B1 (new_n7205_),
	   .A (new_n7204_) );
   INV_X1 g0481 (
	   .ZN (new_n7211_),
	   .A (new_n7210_) );
   BUF_X4 g0480 (
	   .Z (new_n7210_),
	   .A (new_n7209_) );
   NOR2_X1 g0479 (
	   .ZN (new_n7209_),
	   .A2 (new_n7208_),
	   .A1 (new_n7207_1_) );
   INV_X1 g0478 (
	   .ZN (new_n7208_),
	   .A (_net_6006) );
   NOR2_X1 g0477 (
	   .ZN (new_n7207_1_),
	   .A2 (_net_7753),
	   .A1 (new_n7206_) );
   NAND2_X1 g0476 (
	   .ZN (new_n7206_),
	   .A2 (_net_7791),
	   .A1 (net_6059) );
   INV_X1 g0475 (
	   .ZN (new_n7205_),
	   .A (_net_6104) );
   NAND2_X1 g0474 (
	   .ZN (new_n7204_),
	   .A2 (new_n7203_1_),
	   .A1 (new_n7198_) );
   BUF_X4 g0473 (
	   .Z (new_n7203_1_),
	   .A (new_n7202_) );
   NOR2_X1 g0472 (
	   .ZN (new_n7202_),
	   .A2 (new_n7201_),
	   .A1 (new_n7200_) );
   INV_X1 g0471 (
	   .ZN (new_n7201_),
	   .A (_net_6009) );
   NAND4_X1 g0470 (
	   .ZN (new_n7200_),
	   .A4 (_net_7791),
	   .A3 (_net_6006),
	   .A2 (net_6059),
	   .A1 (new_n7199_1_) );
   INV_X1 g0469 (
	   .ZN (new_n7199_1_),
	   .A (_net_7753) );
   NAND2_X1 g0468 (
	   .ZN (new_n7198_),
	   .A2 (new_n7197_),
	   .A1 (new_n7192_) );
   AOI22_X1 g0467 (
	   .ZN (new_n7197_),
	   .B2 (net_6694),
	   .B1 (new_n7196_),
	   .A2 (net_6726),
	   .A1 (new_n7194_1_) );
   BUF_X4 g0466 (
	   .Z (new_n7196_),
	   .A (new_n7195_) );
   NOR2_X1 g0465 (
	   .ZN (new_n7195_),
	   .A2 (_net_6824),
	   .A1 (_net_6823) );
   BUF_X4 g0464 (
	   .Z (new_n7194_1_),
	   .A (new_n7193_) );
   NOR2_X1 g0463 (
	   .ZN (new_n7193_),
	   .A2 (_net_6824),
	   .A1 (new_n7186_) );
   AOI22_X1 g0462 (
	   .ZN (new_n7192_),
	   .B2 (net_6758),
	   .B1 (new_n7191_),
	   .A2 (new_n7189_),
	   .A1 (net_6790) );
   BUF_X4 g0461 (
	   .Z (new_n7191_),
	   .A (new_n7190_1_) );
   NOR2_X1 g0460 (
	   .ZN (new_n7190_1_),
	   .A2 (_net_6823),
	   .A1 (new_n7187_) );
   BUF_X4 g0459 (
	   .Z (new_n7189_),
	   .A (new_n7188_) );
   NOR2_X1 g0458 (
	   .ZN (new_n7188_),
	   .A2 (new_n7187_),
	   .A1 (new_n7186_) );
   INV_X1 g0457 (
	   .ZN (new_n7187_),
	   .A (_net_6824) );
   INV_X1 g0456 (
	   .ZN (new_n7186_),
	   .A (_net_6823) );
   NOR3_X1 g0455 (
	   .ZN (n528),
	   .A3 (new_n7178_),
	   .A2 (new_n7184_),
	   .A1 (new_n7183_) );
   OR4_X1 g0454 (
	   .ZN (new_n7184_),
	   .A4 (x1193),
	   .A3 (x1209),
	   .A2 (new_n7177_1_),
	   .A1 (x1203) );
   INV_X1 g0453 (
	   .ZN (new_n7183_),
	   .A (new_n7182_1_) );
   NAND2_X1 g0452 (
	   .ZN (new_n7182_1_),
	   .A2 (new_n7181_),
	   .A1 (n3157) );
   INV_X1 g0451 (
	   .ZN (new_n7181_),
	   .A (_net_7690) );
   NOR3_X1 g0450 (
	   .ZN (n3157),
	   .A3 (new_n7179_),
	   .A2 (new_n7178_),
	   .A1 (new_n7177_1_) );
   INV_X1 g0449 (
	   .ZN (new_n7179_),
	   .A (_net_7689) );
   INV_X1 g0448 (
	   .ZN (new_n7178_),
	   .A (x1155) );
   NAND2_X1 g0447 (
	   .ZN (new_n7177_1_),
	   .A2 (x1126),
	   .A1 (x1101) );
   NAND3_X1 g0446 (
	   .ZN (n523),
	   .A3 (new_n7175_),
	   .A2 (new_n7160_1_),
	   .A1 (new_n7154_) );
   AND3_X1 g0445 (
	   .ZN (new_n7175_),
	   .A3 (new_n7174_),
	   .A2 (new_n7173_),
	   .A1 (new_n7167_1_) );
   NAND2_X1 g0444 (
	   .ZN (new_n7174_),
	   .A2 (_net_6079),
	   .A1 (new_n6813_1_) );
   NAND2_X1 g0443 (
	   .ZN (new_n7173_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n7172_1_) );
   NAND4_X1 g0442 (
	   .ZN (new_n7172_1_),
	   .A4 (new_n7171_),
	   .A3 (new_n7170_),
	   .A2 (new_n7169_),
	   .A1 (new_n7168_) );
   NAND3_X1 g0441 (
	   .ZN (new_n7171_),
	   .A3 (net_6533),
	   .A2 (_net_6554),
	   .A1 (_net_6553) );
   NAND3_X1 g0440 (
	   .ZN (new_n7170_),
	   .A3 (_net_6554),
	   .A2 (net_6501),
	   .A1 (new_n6789_) );
   NAND3_X1 g0439 (
	   .ZN (new_n7169_),
	   .A3 (net_6469),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   NAND2_X1 g0438 (
	   .ZN (new_n7168_),
	   .A2 (net_6437),
	   .A1 (new_n6785_) );
   NAND2_X1 g0437 (
	   .ZN (new_n7167_1_),
	   .A2 (new_n7166_),
	   .A1 (new_n7165_) );
   BUF_X4 g0436 (
	   .Z (new_n7166_),
	   .A (new_n6809_1_) );
   NAND4_X1 g0435 (
	   .ZN (new_n7165_),
	   .A4 (new_n7164_1_),
	   .A3 (new_n7163_),
	   .A2 (new_n7162_),
	   .A1 (new_n7161_) );
   NAND3_X1 g0434 (
	   .ZN (new_n7164_1_),
	   .A3 (net_6535),
	   .A2 (_net_6554),
	   .A1 (_net_6553) );
   NAND3_X1 g0433 (
	   .ZN (new_n7163_),
	   .A3 (net_6503),
	   .A2 (_net_6554),
	   .A1 (new_n6789_) );
   NAND3_X1 g0432 (
	   .ZN (new_n7162_),
	   .A3 (net_6471),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   NAND2_X1 g0431 (
	   .ZN (new_n7161_),
	   .A2 (net_6439),
	   .A1 (new_n6785_) );
   AOI22_X1 g0430 (
	   .ZN (new_n7160_1_),
	   .B2 (new_n7159_),
	   .B1 (new_n6784_),
	   .A2 (new_n6779_1_),
	   .A1 (net_6547) );
   NAND4_X1 g0429 (
	   .ZN (new_n7159_),
	   .A4 (new_n7158_),
	   .A3 (new_n7157_),
	   .A2 (new_n7156_),
	   .A1 (new_n7155_1_) );
   NAND3_X1 g0428 (
	   .ZN (new_n7158_),
	   .A3 (net_6531),
	   .A2 (_net_6554),
	   .A1 (_net_6553) );
   NAND3_X1 g0427 (
	   .ZN (new_n7157_),
	   .A3 (net_6499),
	   .A2 (_net_6554),
	   .A1 (new_n6789_) );
   NAND3_X1 g0426 (
	   .ZN (new_n7156_),
	   .A3 (net_6467),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   NAND2_X1 g0425 (
	   .ZN (new_n7155_1_),
	   .A2 (net_6435),
	   .A1 (new_n6785_) );
   AND3_X1 g0424 (
	   .ZN (new_n7154_),
	   .A3 (new_n7153_),
	   .A2 (new_n7152_),
	   .A1 (new_n7151_1_) );
   NAND4_X1 g0423 (
	   .ZN (new_n7153_),
	   .A4 (new_n6775_),
	   .A3 (_net_6552),
	   .A2 (net_6515),
	   .A1 (new_n6772_) );
   NAND4_X1 g0422 (
	   .ZN (new_n7152_),
	   .A4 (new_n6770_1_),
	   .A3 (_net_6552),
	   .A2 (net_6451),
	   .A1 (new_n6764_) );
   NAND4_X1 g0421 (
	   .ZN (new_n7151_1_),
	   .A4 (new_n6767_),
	   .A3 (net_6483),
	   .A2 (_net_6552),
	   .A1 (new_n6764_) );
   NOR2_X1 g0420 (
	   .ZN (n518),
	   .A2 (new_n7104_),
	   .A1 (new_n6952_1_) );
   NOR2_X1 g0419 (
	   .ZN (n513),
	   .A2 (new_n6983_),
	   .A1 (new_n7148_) );
   INV_X1 g0418 (
	   .ZN (new_n7148_),
	   .A (_net_5967) );
   CLKBUF_X1 g0417 (
	   .Z (n508),
	   .A (_net_6112) );
   CLKBUF_X1 g0416 (
	   .Z (n503),
	   .A (_net_6091) );
   CLKBUF_X1 g0415 (
	   .Z (n498),
	   .A (net_6059) );
   CLKBUF_X1 g0414 (
	   .Z (n493),
	   .A (_net_7822) );
   CLKBUF_X1 g0413 (
	   .Z (n488),
	   .A (_net_7794) );
   CLKBUF_X1 g0412 (
	   .Z (n484),
	   .A (net_6870) );
   CLKBUF_X1 g0411 (
	   .Z (n479),
	   .A (_net_7818) );
   CLKBUF_X1 g0410 (
	   .Z (n474),
	   .A (net_6397) );
   CLKBUF_X1 g0409 (
	   .Z (n470),
	   .A (net_7388) );
   NAND3_X1 g0408 (
	   .ZN (n465),
	   .A3 (new_n7137_),
	   .A2 (new_n7129_),
	   .A1 (new_n7120_1_) );
   AOI22_X1 g0407 (
	   .ZN (new_n7137_),
	   .B2 (new_n7136_),
	   .B1 (net_6683),
	   .A2 (new_n7134_),
	   .A1 (new_n7013_1_) );
   NOR3_X2 g0406 (
	   .ZN (new_n7136_),
	   .A3 (new_n7135_),
	   .A2 (new_n7113_),
	   .A1 (new_n6977_1_) );
   NAND3_X1 g0405 (
	   .ZN (new_n7135_),
	   .A3 (_net_6689),
	   .A2 (_net_6687),
	   .A1 (_net_6688) );
   NAND4_X1 g0404 (
	   .ZN (new_n7134_),
	   .A4 (new_n7133_1_),
	   .A3 (new_n7132_),
	   .A2 (new_n7131_),
	   .A1 (new_n7130_) );
   NAND3_X1 g0403 (
	   .ZN (new_n7133_1_),
	   .A3 (net_6667),
	   .A2 (_net_6689),
	   .A1 (_net_6688) );
   NAND3_X1 g0402 (
	   .ZN (new_n7132_),
	   .A3 (_net_6689),
	   .A2 (net_6635),
	   .A1 (new_n7004_) );
   NAND3_X1 g0401 (
	   .ZN (new_n7131_),
	   .A3 (_net_6688),
	   .A2 (net_6603),
	   .A1 (new_n7002_) );
   NAND2_X1 g0400 (
	   .ZN (new_n7130_),
	   .A2 (net_6571),
	   .A1 (new_n6973_) );
   AND3_X1 g0399 (
	   .ZN (new_n7129_),
	   .A3 (new_n7128_1_),
	   .A2 (new_n7127_),
	   .A1 (new_n7121_) );
   NAND2_X1 g0398 (
	   .ZN (new_n7128_1_),
	   .A2 (_net_6100),
	   .A1 (new_n6985_) );
   NAND2_X1 g0397 (
	   .ZN (new_n7127_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n7126_) );
   NAND4_X1 g0396 (
	   .ZN (new_n7126_),
	   .A4 (new_n7125_1_),
	   .A3 (new_n7124_),
	   .A2 (new_n7123_),
	   .A1 (new_n7122_) );
   NAND3_X1 g0395 (
	   .ZN (new_n7125_1_),
	   .A3 (net_6669),
	   .A2 (_net_6689),
	   .A1 (_net_6688) );
   NAND3_X1 g0394 (
	   .ZN (new_n7124_),
	   .A3 (_net_6689),
	   .A2 (net_6637),
	   .A1 (new_n7004_) );
   NAND3_X1 g0393 (
	   .ZN (new_n7123_),
	   .A3 (net_6605),
	   .A2 (_net_6688),
	   .A1 (new_n7002_) );
   NAND2_X1 g0392 (
	   .ZN (new_n7122_),
	   .A2 (net_6573),
	   .A1 (new_n6973_) );
   NAND2_X1 g0391 (
	   .ZN (new_n7121_),
	   .A2 (new_n6980_),
	   .A1 (new_n7007_) );
   AND3_X1 g0390 (
	   .ZN (new_n7120_1_),
	   .A3 (new_n7119_),
	   .A2 (new_n7117_),
	   .A1 (new_n7116_1_) );
   NAND4_X1 g0389 (
	   .ZN (new_n7119_),
	   .A4 (new_n6987_),
	   .A3 (net_6651),
	   .A2 (_net_6687),
	   .A1 (new_n7118_) );
   BUF_X4 g0388 (
	   .Z (new_n7118_),
	   .A (new_n7114_) );
   NAND4_X1 g0387 (
	   .ZN (new_n7117_),
	   .A4 (new_n6990_1_),
	   .A3 (net_6587),
	   .A2 (_net_6687),
	   .A1 (new_n7115_) );
   NAND4_X1 g0386 (
	   .ZN (new_n7116_1_),
	   .A4 (new_n6989_),
	   .A3 (_net_6687),
	   .A2 (net_6619),
	   .A1 (new_n7115_) );
   BUF_X4 g0385 (
	   .Z (new_n7115_),
	   .A (new_n7114_) );
   NOR2_X1 g0384 (
	   .ZN (new_n7114_),
	   .A2 (new_n7113_),
	   .A1 (new_n6977_1_) );
   INV_X1 g0383 (
	   .ZN (new_n7113_),
	   .A (new_n6997_) );
   OAI21_X1 g0382 (
	   .ZN (n460),
	   .B2 (new_n7111_1_),
	   .B1 (new_n7110_),
	   .A (new_n7109_) );
   BUF_X4 g0381 (
	   .Z (new_n7111_1_),
	   .A (new_n7100_) );
   INV_X1 g0380 (
	   .ZN (new_n7110_),
	   .A (_net_7355) );
   NAND2_X1 g0379 (
	   .ZN (new_n7109_),
	   .A2 (new_n7108_),
	   .A1 (new_n7101_) );
   OAI221_X1 g0378 (
	   .ZN (new_n7108_),
	   .C2 (new_n7107_1_),
	   .C1 (new_n7106_),
	   .B2 (new_n7105_),
	   .B1 (new_n7104_),
	   .A (new_n7103_) );
   INV_X1 g0377 (
	   .ZN (new_n7107_1_),
	   .A (net_335) );
   INV_X2 g0376 (
	   .ZN (new_n7106_),
	   .A (_net_270) );
   INV_X1 g0375 (
	   .ZN (new_n7105_),
	   .A (_net_269) );
   INV_X1 g0374 (
	   .ZN (new_n7104_),
	   .A (net_337) );
   NAND2_X1 g0373 (
	   .ZN (new_n7103_),
	   .A2 (net_7243),
	   .A1 (new_n7102_1_) );
   BUF_X4 g0372 (
	   .Z (new_n7102_1_),
	   .A (new_n6942_) );
   BUF_X4 g0371 (
	   .Z (new_n7101_),
	   .A (new_n7100_) );
   BUF_X4 g0370 (
	   .Z (new_n7100_),
	   .A (new_n7099_) );
   AND2_X1 g0369 (
	   .ZN (new_n7099_),
	   .A2 (new_n7098_1_),
	   .A1 (new_n6945_) );
   INV_X1 g0368 (
	   .ZN (new_n7098_1_),
	   .A (new_n7097_) );
   NAND2_X1 g0367 (
	   .ZN (new_n7097_),
	   .A2 (_net_7383),
	   .A1 (_net_7382) );
   CLKBUF_X1 g0366 (
	   .Z (n455),
	   .A (_net_7798) );
   CLKBUF_X1 g0365 (
	   .Z (n451),
	   .A (x1527) );
   NAND4_X1 g0364 (
	   .ZN (n447),
	   .A4 (new_n7093_1_),
	   .A3 (new_n7081_),
	   .A2 (new_n7071_),
	   .A1 (new_n7061_) );
   AOI22_X1 g0363 (
	   .ZN (new_n7093_1_),
	   .B2 (_net_6150),
	   .B1 (new_n7092_),
	   .A2 (new_n7089_1_),
	   .A1 (new_n7086_) );
   BUF_X4 g0362 (
	   .Z (new_n7092_),
	   .A (new_n7091_) );
   NOR2_X1 g0361 (
	   .ZN (new_n7091_),
	   .A2 (new_n7090_),
	   .A1 (new_n7056_) );
   INV_X1 g0360 (
	   .ZN (new_n7090_),
	   .A (_net_6028) );
   BUF_X4 g0359 (
	   .Z (new_n7089_1_),
	   .A (new_n7088_) );
   NOR2_X1 g0358 (
	   .ZN (new_n7088_),
	   .A2 (new_n7087_),
	   .A1 (new_n7067_1_) );
   INV_X1 g0357 (
	   .ZN (new_n7087_),
	   .A (_net_6031) );
   NAND4_X1 g0356 (
	   .ZN (new_n7086_),
	   .A4 (new_n7085_1_),
	   .A3 (new_n7084_),
	   .A2 (new_n7083_),
	   .A1 (new_n7082_1_) );
   NAND3_X1 g0355 (
	   .ZN (new_n7085_1_),
	   .A3 (_net_7093),
	   .A2 (net_7066),
	   .A1 (_net_7094) );
   NAND3_X1 g0354 (
	   .ZN (new_n7084_),
	   .A3 (net_7034),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   NAND3_X1 g0353 (
	   .ZN (new_n7083_),
	   .A3 (net_7002),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   NAND2_X1 g0352 (
	   .ZN (new_n7082_1_),
	   .A2 (net_6970),
	   .A1 (new_n7063_) );
   NAND2_X1 g0351 (
	   .ZN (new_n7081_),
	   .A2 (new_n7080_),
	   .A1 (new_n7073_) );
   NAND4_X1 g0350 (
	   .ZN (new_n7080_),
	   .A4 (new_n7079_),
	   .A3 (new_n7078_),
	   .A2 (new_n7076_),
	   .A1 (new_n7074_) );
   NAND3_X1 g0349 (
	   .ZN (new_n7079_),
	   .A3 (net_7078),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   NAND3_X1 g0348 (
	   .ZN (new_n7078_),
	   .A3 (net_7046),
	   .A2 (_net_7094),
	   .A1 (new_n7077_1_) );
   BUF_X4 g0347 (
	   .Z (new_n7077_1_),
	   .A (new_n7048_) );
   NAND3_X1 g0346 (
	   .ZN (new_n7076_),
	   .A3 (net_7014),
	   .A2 (_net_7093),
	   .A1 (new_n7075_) );
   BUF_X4 g0345 (
	   .Z (new_n7075_),
	   .A (new_n7042_) );
   NAND2_X1 g0344 (
	   .ZN (new_n7074_),
	   .A2 (net_6982),
	   .A1 (new_n7063_) );
   NOR2_X1 g0343 (
	   .ZN (new_n7073_),
	   .A2 (new_n7072_1_),
	   .A1 (new_n7058_1_) );
   INV_X1 g0342 (
	   .ZN (new_n7072_1_),
	   .A (_net_7092) );
   NAND2_X1 g0341 (
	   .ZN (new_n7071_),
	   .A2 (new_n7070_),
	   .A1 (new_n7065_) );
   BUF_X4 g0340 (
	   .Z (new_n7070_),
	   .A (new_n7069_) );
   NOR2_X1 g0339 (
	   .ZN (new_n7069_),
	   .A2 (new_n7068_),
	   .A1 (new_n7067_1_) );
   INV_X1 g0338 (
	   .ZN (new_n7068_),
	   .A (_net_6030) );
   NAND4_X1 g0337 (
	   .ZN (new_n7067_1_),
	   .A4 (_net_6028),
	   .A3 (_net_7791),
	   .A2 (net_6057),
	   .A1 (new_n7066_) );
   INV_X1 g0336 (
	   .ZN (new_n7066_),
	   .A (_net_7757) );
   NAND2_X1 g0335 (
	   .ZN (new_n7065_),
	   .A2 (new_n7064_),
	   .A1 (new_n7062_1_) );
   AOI22_X1 g0334 (
	   .ZN (new_n7064_),
	   .B2 (net_6968),
	   .B1 (new_n7063_),
	   .A2 (net_7000),
	   .A1 (new_n7049_1_) );
   BUF_X4 g0333 (
	   .Z (new_n7063_),
	   .A (new_n7051_) );
   AOI22_X1 g0332 (
	   .ZN (new_n7062_1_),
	   .B2 (net_7064),
	   .B1 (new_n7046_),
	   .A2 (new_n7043_),
	   .A1 (net_7032) );
   NAND2_X1 g0331 (
	   .ZN (new_n7061_),
	   .A2 (new_n7060_),
	   .A1 (new_n7054_) );
   BUF_X4 g0330 (
	   .Z (new_n7060_),
	   .A (new_n7059_) );
   NOR2_X1 g0329 (
	   .ZN (new_n7059_),
	   .A2 (_net_7092),
	   .A1 (new_n7058_1_) );
   NAND3_X1 g0328 (
	   .ZN (new_n7058_1_),
	   .A3 (new_n7057_),
	   .A2 (_net_6028),
	   .A1 (new_n7056_) );
   NOR2_X1 g0327 (
	   .ZN (new_n7057_),
	   .A2 (_net_6031),
	   .A1 (_net_6030) );
   NOR2_X1 g0326 (
	   .ZN (new_n7056_),
	   .A2 (_net_7757),
	   .A1 (new_n7055_) );
   NAND2_X1 g0325 (
	   .ZN (new_n7055_),
	   .A2 (_net_7791),
	   .A1 (net_6057) );
   NAND2_X1 g0324 (
	   .ZN (new_n7054_),
	   .A2 (new_n7053_1_),
	   .A1 (new_n7047_) );
   AOI22_X1 g0323 (
	   .ZN (new_n7053_1_),
	   .B2 (net_6966),
	   .B1 (new_n7052_),
	   .A2 (net_6998),
	   .A1 (new_n7050_) );
   BUF_X4 g0322 (
	   .Z (new_n7052_),
	   .A (new_n7051_) );
   NOR2_X1 g0321 (
	   .ZN (new_n7051_),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   BUF_X4 g0320 (
	   .Z (new_n7050_),
	   .A (new_n7049_1_) );
   NOR2_X1 g0319 (
	   .ZN (new_n7049_1_),
	   .A2 (_net_7094),
	   .A1 (new_n7048_) );
   INV_X1 g0318 (
	   .ZN (new_n7048_),
	   .A (_net_7093) );
   AOI22_X1 g0317 (
	   .ZN (new_n7047_),
	   .B2 (net_7062),
	   .B1 (new_n7046_),
	   .A2 (new_n7044_),
	   .A1 (net_7030) );
   INV_X1 g0316 (
	   .ZN (new_n7046_),
	   .A (new_n7045_1_) );
   NAND2_X1 g0315 (
	   .ZN (new_n7045_1_),
	   .A2 (_net_7093),
	   .A1 (_net_7094) );
   BUF_X4 g0314 (
	   .Z (new_n7044_),
	   .A (new_n7043_) );
   NOR2_X1 g0313 (
	   .ZN (new_n7043_),
	   .A2 (_net_7093),
	   .A1 (new_n7042_) );
   INV_X1 g0312 (
	   .ZN (new_n7042_),
	   .A (_net_7094) );
   CLKBUF_X1 g0311 (
	   .Z (n443),
	   .A (net_7000) );
   CLKBUF_X1 g0310 (
	   .Z (n438),
	   .A (_net_7815) );
   CLKBUF_X1 g0309 (
	   .Z (n434),
	   .A (net_7713) );
   CLKBUF_X1 g0308 (
	   .Z (n429),
	   .A (_net_7806) );
   CLKBUF_X1 g0307 (
	   .Z (n424),
	   .A (_net_7819) );
   NOR2_X1 g0306 (
	   .ZN (n420),
	   .A2 (new_n6900_),
	   .A1 (new_n7035_) );
   BUF_X4 g0305 (
	   .Z (new_n7035_),
	   .A (new_n7034_) );
   INV_X2 g0304 (
	   .ZN (new_n7034_),
	   .A (new_n6889_) );
   CLKBUF_X1 g0303 (
	   .Z (n415),
	   .A (_net_7795) );
   CLKBUF_X1 g0302 (
	   .Z (n410),
	   .A (_net_6117) );
   CLKBUF_X1 g0301 (
	   .Z (n405),
	   .A (net_6395) );
   MUX2_X1 g0300 (
	   .Z (n400),
	   .S (new_n7029_),
	   .B (_net_7595),
	   .A (new_n7022_) );
   BUF_X8 g0299 (
	   .Z (new_n7029_),
	   .A (new_n7028_) );
   NAND3_X1 g0298 (
	   .ZN (new_n7028_),
	   .A3 (new_n7027_1_),
	   .A2 (_net_7684),
	   .A1 (new_n7026_) );
   INV_X1 g0297 (
	   .ZN (new_n7027_1_),
	   .A (_net_7685) );
   AOI21_X1 g0296 (
	   .ZN (new_n7026_),
	   .B2 (new_n7018_1_),
	   .B1 (new_n7025_),
	   .A (new_n7024_) );
   INV_X1 g0295 (
	   .ZN (new_n7025_),
	   .A (_net_7683) );
   NAND3_X1 g0294 (
	   .ZN (new_n7024_),
	   .A3 (_net_5924),
	   .A2 (net_5858),
	   .A1 (new_n7023_1_) );
   INV_X1 g0293 (
	   .ZN (new_n7023_1_),
	   .A (_net_7765) );
   OAI21_X1 g0292 (
	   .ZN (new_n7022_),
	   .B2 (new_n7021_),
	   .B1 (new_n7020_),
	   .A (new_n7017_) );
   INV_X1 g0291 (
	   .ZN (new_n7021_),
	   .A (net_7547) );
   BUF_X4 g0290 (
	   .Z (new_n7020_),
	   .A (new_n7019_) );
   INV_X2 g0289 (
	   .ZN (new_n7019_),
	   .A (new_n7018_1_) );
   NOR2_X1 g0288 (
	   .ZN (new_n7018_1_),
	   .A2 (_net_292),
	   .A1 (_net_291) );
   AOI22_X1 g0287 (
	   .ZN (new_n7017_),
	   .B2 (_net_291),
	   .B1 (net_379),
	   .A2 (_net_292),
	   .A1 (net_377) );
   CLKBUF_X1 g0286 (
	   .Z (n395),
	   .A (_net_7820) );
   NAND4_X1 g0285 (
	   .ZN (n390),
	   .A4 (new_n7014_),
	   .A3 (new_n7008_),
	   .A2 (new_n6996_),
	   .A1 (new_n6986_1_) );
   NAND2_X1 g0284 (
	   .ZN (new_n7014_),
	   .A2 (new_n7013_1_),
	   .A1 (new_n7011_) );
   BUF_X4 g0283 (
	   .Z (new_n7013_1_),
	   .A (new_n7012_) );
   NOR2_X1 g0282 (
	   .ZN (new_n7012_),
	   .A2 (_net_6687),
	   .A1 (new_n6998_) );
   NAND2_X1 g0281 (
	   .ZN (new_n7011_),
	   .A2 (new_n7010_),
	   .A1 (new_n7009_1_) );
   AOI22_X1 g0280 (
	   .ZN (new_n7010_),
	   .B2 (net_6559),
	   .B1 (new_n6990_1_),
	   .A2 (net_6591),
	   .A1 (new_n6989_) );
   AOI22_X1 g0279 (
	   .ZN (new_n7009_1_),
	   .B2 (net_6655),
	   .B1 (new_n6968_),
	   .A2 (new_n6987_),
	   .A1 (net_6623) );
   NAND2_X1 g0278 (
	   .ZN (new_n7008_),
	   .A2 (new_n7007_),
	   .A1 (new_n7000_1_) );
   NAND4_X1 g0277 (
	   .ZN (new_n7007_),
	   .A4 (new_n7006_),
	   .A3 (new_n7005_1_),
	   .A2 (new_n7003_),
	   .A1 (new_n7001_) );
   NAND3_X1 g0276 (
	   .ZN (new_n7006_),
	   .A3 (_net_6689),
	   .A2 (_net_6688),
	   .A1 (net_6671) );
   NAND3_X1 g0275 (
	   .ZN (new_n7005_1_),
	   .A3 (_net_6689),
	   .A2 (net_6639),
	   .A1 (new_n7004_) );
   BUF_X4 g0274 (
	   .Z (new_n7004_),
	   .A (new_n6970_) );
   NAND3_X1 g0273 (
	   .ZN (new_n7003_),
	   .A3 (net_6607),
	   .A2 (_net_6688),
	   .A1 (new_n7002_) );
   BUF_X4 g0272 (
	   .Z (new_n7002_),
	   .A (new_n6965_) );
   NAND2_X1 g0271 (
	   .ZN (new_n7001_),
	   .A2 (net_6575),
	   .A1 (new_n6973_) );
   NOR2_X1 g0270 (
	   .ZN (new_n7000_1_),
	   .A2 (new_n6999_),
	   .A1 (new_n6998_) );
   INV_X1 g0269 (
	   .ZN (new_n6999_),
	   .A (_net_6687) );
   NAND3_X1 g0268 (
	   .ZN (new_n6998_),
	   .A3 (new_n6997_),
	   .A2 (_net_5995),
	   .A1 (new_n6982_1_) );
   NOR2_X1 g0267 (
	   .ZN (new_n6997_),
	   .A2 (_net_5998),
	   .A1 (_net_5997) );
   NAND2_X1 g0266 (
	   .ZN (new_n6996_),
	   .A2 (new_n6995_1_),
	   .A1 (new_n6992_) );
   BUF_X4 g0265 (
	   .Z (new_n6995_1_),
	   .A (new_n6994_) );
   NOR2_X1 g0264 (
	   .ZN (new_n6994_),
	   .A2 (new_n6993_),
	   .A1 (new_n6977_1_) );
   INV_X1 g0263 (
	   .ZN (new_n6993_),
	   .A (_net_5997) );
   NAND2_X1 g0262 (
	   .ZN (new_n6992_),
	   .A2 (new_n6991_),
	   .A1 (new_n6988_) );
   AOI22_X1 g0261 (
	   .ZN (new_n6991_),
	   .B2 (net_6561),
	   .B1 (new_n6990_1_),
	   .A2 (net_6593),
	   .A1 (new_n6989_) );
   BUF_X4 g0260 (
	   .Z (new_n6990_1_),
	   .A (new_n6972_) );
   BUF_X4 g0259 (
	   .Z (new_n6989_),
	   .A (new_n6971_) );
   AOI22_X1 g0258 (
	   .ZN (new_n6988_),
	   .B2 (net_6657),
	   .B1 (new_n6968_),
	   .A2 (new_n6987_),
	   .A1 (net_6625) );
   BUF_X4 g0257 (
	   .Z (new_n6987_),
	   .A (new_n6966_) );
   AOI22_X1 g0256 (
	   .ZN (new_n6986_1_),
	   .B2 (new_n6985_),
	   .B1 (_net_6088),
	   .A2 (new_n6980_),
	   .A1 (new_n6975_) );
   BUF_X4 g0255 (
	   .Z (new_n6985_),
	   .A (new_n6984_) );
   NOR2_X1 g0254 (
	   .ZN (new_n6984_),
	   .A2 (new_n6983_),
	   .A1 (new_n6982_1_) );
   INV_X1 g0253 (
	   .ZN (new_n6983_),
	   .A (_net_5995) );
   NOR2_X1 g0252 (
	   .ZN (new_n6982_1_),
	   .A2 (_net_7751),
	   .A1 (new_n6981_) );
   NAND2_X1 g0251 (
	   .ZN (new_n6981_),
	   .A2 (_net_7791),
	   .A1 (net_6060) );
   BUF_X4 g0250 (
	   .Z (new_n6980_),
	   .A (new_n6979_) );
   NOR2_X1 g0249 (
	   .ZN (new_n6979_),
	   .A2 (new_n6978_),
	   .A1 (new_n6977_1_) );
   INV_X1 g0248 (
	   .ZN (new_n6978_),
	   .A (_net_5998) );
   NAND4_X1 g0247 (
	   .ZN (new_n6977_1_),
	   .A4 (_net_5995),
	   .A3 (_net_7791),
	   .A2 (net_6060),
	   .A1 (new_n6976_) );
   INV_X1 g0246 (
	   .ZN (new_n6976_),
	   .A (_net_7751) );
   NAND2_X1 g0245 (
	   .ZN (new_n6975_),
	   .A2 (new_n6974_1_),
	   .A1 (new_n6969_1_) );
   AOI22_X1 g0244 (
	   .ZN (new_n6974_1_),
	   .B2 (net_6563),
	   .B1 (new_n6973_),
	   .A2 (net_6595),
	   .A1 (new_n6971_) );
   BUF_X4 g0243 (
	   .Z (new_n6973_),
	   .A (new_n6972_) );
   NOR2_X1 g0242 (
	   .ZN (new_n6972_),
	   .A2 (_net_6689),
	   .A1 (_net_6688) );
   NOR2_X1 g0241 (
	   .ZN (new_n6971_),
	   .A2 (_net_6689),
	   .A1 (new_n6970_) );
   INV_X1 g0240 (
	   .ZN (new_n6970_),
	   .A (_net_6688) );
   AOI22_X1 g0239 (
	   .ZN (new_n6969_1_),
	   .B2 (net_6659),
	   .B1 (new_n6968_),
	   .A2 (new_n6966_),
	   .A1 (net_6627) );
   INV_X1 g0238 (
	   .ZN (new_n6968_),
	   .A (new_n6967_) );
   NAND2_X1 g0237 (
	   .ZN (new_n6967_),
	   .A2 (_net_6689),
	   .A1 (_net_6688) );
   NOR2_X1 g0236 (
	   .ZN (new_n6966_),
	   .A2 (_net_6688),
	   .A1 (new_n6965_) );
   INV_X1 g0235 (
	   .ZN (new_n6965_),
	   .A (_net_6689) );
   NAND2_X1 g0234 (
	   .ZN (n385),
	   .A2 (_net_6404),
	   .A1 (new_n6963_) );
   INV_X1 g0233 (
	   .ZN (new_n6963_),
	   .A (x38) );
   OAI21_X1 g0232 (
	   .ZN (n380),
	   .B2 (new_n6961_),
	   .B1 (new_n6960_1_),
	   .A (new_n6959_) );
   INV_X1 g0231 (
	   .ZN (new_n6961_),
	   .A (_net_262) );
   INV_X1 g0230 (
	   .ZN (new_n6960_1_),
	   .A (_net_264) );
   INV_X1 g0229 (
	   .ZN (new_n6959_),
	   .A (_net_298) );
   OAI21_X1 g0228 (
	   .ZN (n375),
	   .B2 (new_n6957_1_),
	   .B1 (new_n6956_),
	   .A (new_n6955_) );
   BUF_X4 g0227 (
	   .Z (new_n6957_1_),
	   .A (new_n6948_) );
   INV_X1 g0226 (
	   .ZN (new_n6956_),
	   .A (_net_7252) );
   NAND2_X1 g0225 (
	   .ZN (new_n6955_),
	   .A2 (new_n6954_),
	   .A1 (new_n6949_) );
   OAI21_X1 g0224 (
	   .ZN (new_n6954_),
	   .B2 (new_n6953_),
	   .B1 (new_n6952_1_),
	   .A (new_n6950_) );
   INV_X1 g0223 (
	   .ZN (new_n6953_),
	   .A (net_7236) );
   BUF_X4 g0222 (
	   .Z (new_n6952_1_),
	   .A (new_n6951_) );
   INV_X1 g0221 (
	   .ZN (new_n6951_),
	   .A (new_n6942_) );
   AOI22_X1 g0220 (
	   .ZN (new_n6950_),
	   .B2 (net_330),
	   .B1 (_net_269),
	   .A2 (net_328),
	   .A1 (_net_270) );
   BUF_X4 g0219 (
	   .Z (new_n6949_),
	   .A (new_n6948_) );
   BUF_X4 g0218 (
	   .Z (new_n6948_),
	   .A (new_n6947_1_) );
   AND2_X1 g0217 (
	   .ZN (new_n6947_1_),
	   .A2 (new_n6946_),
	   .A1 (new_n6945_) );
   NOR2_X1 g0216 (
	   .ZN (new_n6946_),
	   .A2 (_net_7383),
	   .A1 (_net_7382) );
   AND2_X2 g0215 (
	   .ZN (new_n6945_),
	   .A2 (new_n6944_),
	   .A1 (new_n6941_) );
   NAND2_X1 g0214 (
	   .ZN (new_n6944_),
	   .A2 (new_n6943_1_),
	   .A1 (new_n6942_) );
   INV_X1 g0213 (
	   .ZN (new_n6943_1_),
	   .A (_net_7381) );
   NOR2_X2 g0212 (
	   .ZN (new_n6942_),
	   .A2 (_net_269),
	   .A1 (_net_270) );
   NOR3_X1 g0211 (
	   .ZN (new_n6941_),
	   .A3 (_net_7761),
	   .A2 (new_n6940_),
	   .A1 (new_n6939_) );
   INV_X1 g0210 (
	   .ZN (new_n6940_),
	   .A (_net_5922) );
   INV_X1 g0209 (
	   .ZN (new_n6939_),
	   .A (net_5861) );
   OAI21_X1 g0208 (
	   .ZN (n370),
	   .B2 (new_n6907_),
	   .B1 (new_n6937_),
	   .A (new_n6936_) );
   INV_X1 g0207 (
	   .ZN (new_n6937_),
	   .A (_net_7474) );
   NAND2_X1 g0206 (
	   .ZN (new_n6936_),
	   .A2 (new_n6935_),
	   .A1 (new_n6897_) );
   OAI221_X1 g0205 (
	   .ZN (new_n6935_),
	   .C2 (new_n6901_),
	   .C1 (new_n6934_1_),
	   .B2 (new_n6902_1_),
	   .B1 (new_n6933_),
	   .A (new_n6932_) );
   INV_X1 g0204 (
	   .ZN (new_n6934_1_),
	   .A (net_355) );
   INV_X1 g0203 (
	   .ZN (new_n6933_),
	   .A (net_357) );
   NAND2_X1 g0202 (
	   .ZN (new_n6932_),
	   .A2 (net_7394),
	   .A1 (new_n6898_) );
   CLKBUF_X1 g0201 (
	   .Z (n366),
	   .A (net_6996) );
   CLKBUF_X1 g0200 (
	   .Z (n361),
	   .A (_net_7819) );
   CLKBUF_X1 g0199 (
	   .Z (n357),
	   .A (net_7114) );
   CLKBUF_X1 g0198 (
	   .Z (n352),
	   .A (x1542) );
   CLKBUF_X1 g0197 (
	   .Z (n349),
	   .A (net_6474) );
   CLKBUF_X1 g0196 (
	   .Z (n344),
	   .A (_net_6080) );
   CLKBUF_X1 g0195 (
	   .Z (n339),
	   .A (_net_6168) );
   CLKBUF_X1 g0194 (
	   .Z (n334),
	   .A (net_133) );
   MUX2_X1 g0193 (
	   .Z (n329),
	   .S (_net_7791),
	   .B (net_155),
	   .A (_net_6062) );
   CLKBUF_X1 g0192 (
	   .Z (n324),
	   .A (net_7802) );
   OAI221_X1 g0191 (
	   .ZN (n319),
	   .C2 (new_n6920_),
	   .C1 (new_n6918_),
	   .B2 (new_n6917_),
	   .B1 (new_n6915_1_),
	   .A (new_n6914_) );
   BUF_X4 g0190 (
	   .Z (new_n6920_),
	   .A (new_n6919_1_) );
   NAND2_X1 g0189 (
	   .ZN (new_n6919_1_),
	   .A2 (net_7378),
	   .A1 (_net_7379) );
   INV_X1 g0188 (
	   .ZN (new_n6918_),
	   .A (_net_7365) );
   BUF_X4 g0187 (
	   .Z (new_n6917_),
	   .A (new_n6916_) );
   NAND2_X1 g0186 (
	   .ZN (new_n6916_),
	   .A2 (net_7378),
	   .A1 (new_n6909_) );
   INV_X1 g0185 (
	   .ZN (new_n6915_1_),
	   .A (_net_7301) );
   AOI22_X1 g0184 (
	   .ZN (new_n6914_),
	   .B2 (_net_7269),
	   .B1 (new_n6913_),
	   .A2 (_net_7333),
	   .A1 (new_n6911_) );
   BUF_X4 g0183 (
	   .Z (new_n6913_),
	   .A (new_n6912_) );
   NOR2_X1 g0182 (
	   .ZN (new_n6912_),
	   .A2 (net_7378),
	   .A1 (_net_7379) );
   BUF_X4 g0181 (
	   .Z (new_n6911_),
	   .A (new_n6910_1_) );
   NOR2_X1 g0180 (
	   .ZN (new_n6910_1_),
	   .A2 (net_7378),
	   .A1 (new_n6909_) );
   INV_X1 g0179 (
	   .ZN (new_n6909_),
	   .A (_net_7379) );
   OAI21_X1 g0178 (
	   .ZN (n314),
	   .B2 (new_n6907_),
	   .B1 (new_n6906_1_),
	   .A (new_n6905_) );
   BUF_X4 g0177 (
	   .Z (new_n6907_),
	   .A (new_n6896_) );
   INV_X1 g0176 (
	   .ZN (new_n6906_1_),
	   .A (_net_7481) );
   NAND2_X1 g0175 (
	   .ZN (new_n6905_),
	   .A2 (new_n6904_),
	   .A1 (new_n6897_) );
   OAI221_X1 g0174 (
	   .ZN (new_n6904_),
	   .C2 (new_n6903_),
	   .C1 (new_n6902_1_),
	   .B2 (new_n6901_),
	   .B1 (new_n6900_),
	   .A (new_n6899_1_) );
   INV_X1 g0173 (
	   .ZN (new_n6903_),
	   .A (net_364) );
   INV_X2 g0172 (
	   .ZN (new_n6902_1_),
	   .A (_net_280) );
   INV_X2 g0171 (
	   .ZN (new_n6901_),
	   .A (_net_281) );
   INV_X1 g0170 (
	   .ZN (new_n6900_),
	   .A (net_362) );
   NAND2_X1 g0169 (
	   .ZN (new_n6899_1_),
	   .A2 (net_350),
	   .A1 (new_n6898_) );
   BUF_X4 g0168 (
	   .Z (new_n6898_),
	   .A (new_n6889_) );
   BUF_X4 g0167 (
	   .Z (new_n6897_),
	   .A (new_n6896_) );
   BUF_X4 g0166 (
	   .Z (new_n6896_),
	   .A (new_n6895_1_) );
   AND2_X1 g0165 (
	   .ZN (new_n6895_1_),
	   .A2 (new_n6894_),
	   .A1 (new_n6892_) );
   NOR2_X1 g0164 (
	   .ZN (new_n6894_),
	   .A2 (_net_7533),
	   .A1 (new_n6893_) );
   INV_X1 g0163 (
	   .ZN (new_n6893_),
	   .A (_net_7534) );
   AND2_X2 g0162 (
	   .ZN (new_n6892_),
	   .A2 (new_n6891_),
	   .A1 (new_n6888_) );
   NAND2_X1 g0161 (
	   .ZN (new_n6891_),
	   .A2 (new_n6890_1_),
	   .A1 (new_n6889_) );
   INV_X1 g0160 (
	   .ZN (new_n6890_1_),
	   .A (_net_7532) );
   NOR2_X1 g0159 (
	   .ZN (new_n6889_),
	   .A2 (_net_281),
	   .A1 (_net_280) );
   NOR3_X1 g0158 (
	   .ZN (new_n6888_),
	   .A3 (_net_7763),
	   .A2 (new_n6887_),
	   .A1 (new_n6886_1_) );
   INV_X1 g0157 (
	   .ZN (new_n6887_),
	   .A (net_5860) );
   INV_X1 g0156 (
	   .ZN (new_n6886_1_),
	   .A (_net_5920) );
   CLKBUF_X1 g0155 (
	   .Z (n310),
	   .A (net_6704) );
   CLKBUF_X1 g0154 (
	   .Z (n305),
	   .A (_net_7820) );
   NAND3_X1 g0153 (
	   .ZN (n300),
	   .A3 (new_n6882_),
	   .A2 (new_n6871_),
	   .A1 (new_n6843_) );
   AOI22_X1 g0152 (
	   .ZN (new_n6882_),
	   .B2 (new_n6881_1_),
	   .B1 (net_6946),
	   .A2 (new_n6879_),
	   .A1 (new_n6876_1_) );
   NOR3_X2 g0151 (
	   .ZN (new_n6881_1_),
	   .A3 (new_n6880_),
	   .A2 (new_n6828_),
	   .A1 (new_n6826_1_) );
   NAND3_X1 g0150 (
	   .ZN (new_n6880_),
	   .A3 (_net_6958),
	   .A2 (_net_6959),
	   .A1 (_net_6957) );
   BUF_X4 g0149 (
	   .Z (new_n6879_),
	   .A (new_n6878_) );
   NOR2_X1 g0148 (
	   .ZN (new_n6878_),
	   .A2 (_net_6957),
	   .A1 (new_n6877_) );
   NAND3_X1 g0147 (
	   .ZN (new_n6877_),
	   .A3 (new_n6827_),
	   .A2 (_net_6017),
	   .A1 (new_n6866_) );
   NAND2_X1 g0146 (
	   .ZN (new_n6876_1_),
	   .A2 (new_n6875_),
	   .A1 (new_n6874_) );
   AOI22_X1 g0145 (
	   .ZN (new_n6875_),
	   .B2 (net_6834),
	   .B1 (new_n6844_),
	   .A2 (net_6866),
	   .A1 (new_n6832_) );
   AOI22_X1 g0144 (
	   .ZN (new_n6874_),
	   .B2 (net_6930),
	   .B1 (new_n6873_),
	   .A2 (new_n6840_1_),
	   .A1 (net_6898) );
   INV_X1 g0143 (
	   .ZN (new_n6873_),
	   .A (new_n6872_1_) );
   NAND2_X1 g0142 (
	   .ZN (new_n6872_1_),
	   .A2 (_net_6958),
	   .A1 (_net_6959) );
   AND3_X1 g0141 (
	   .ZN (new_n6871_),
	   .A3 (new_n6870_),
	   .A2 (new_n6864_),
	   .A1 (new_n6855_1_) );
   NAND2_X1 g0140 (
	   .ZN (new_n6870_),
	   .A2 (_net_6133),
	   .A1 (new_n6869_) );
   BUF_X4 g0139 (
	   .Z (new_n6869_),
	   .A (new_n6868_) );
   NOR2_X1 g0138 (
	   .ZN (new_n6868_),
	   .A2 (new_n6867_1_),
	   .A1 (new_n6866_) );
   INV_X1 g0137 (
	   .ZN (new_n6867_1_),
	   .A (_net_6017) );
   NOR2_X1 g0136 (
	   .ZN (new_n6866_),
	   .A2 (_net_7755),
	   .A1 (new_n6865_) );
   NAND2_X1 g0135 (
	   .ZN (new_n6865_),
	   .A2 (net_6058),
	   .A1 (_net_7791) );
   NAND2_X1 g0134 (
	   .ZN (new_n6864_),
	   .A2 (new_n6863_1_),
	   .A1 (new_n6860_1_) );
   BUF_X4 g0133 (
	   .Z (new_n6863_1_),
	   .A (new_n6862_) );
   NOR2_X1 g0132 (
	   .ZN (new_n6862_),
	   .A2 (new_n6861_),
	   .A1 (new_n6826_1_) );
   INV_X1 g0131 (
	   .ZN (new_n6861_),
	   .A (_net_6019) );
   NAND4_X1 g0130 (
	   .ZN (new_n6860_1_),
	   .A4 (new_n6859_),
	   .A3 (new_n6858_),
	   .A2 (new_n6857_),
	   .A1 (new_n6856_) );
   NAND3_X1 g0129 (
	   .ZN (new_n6859_),
	   .A3 (net_6932),
	   .A2 (_net_6958),
	   .A1 (_net_6959) );
   NAND3_X1 g0128 (
	   .ZN (new_n6858_),
	   .A3 (_net_6959),
	   .A2 (net_6900),
	   .A1 (new_n6848_) );
   NAND3_X1 g0127 (
	   .ZN (new_n6857_),
	   .A3 (_net_6958),
	   .A2 (net_6868),
	   .A1 (new_n6846_) );
   NAND2_X1 g0126 (
	   .ZN (new_n6856_),
	   .A2 (net_6836),
	   .A1 (new_n6844_) );
   NAND2_X1 g0125 (
	   .ZN (new_n6855_1_),
	   .A2 (new_n6854_),
	   .A1 (new_n6851_) );
   BUF_X4 g0124 (
	   .Z (new_n6854_),
	   .A (new_n6853_) );
   NOR2_X1 g0123 (
	   .ZN (new_n6853_),
	   .A2 (new_n6852_),
	   .A1 (new_n6826_1_) );
   INV_X1 g0122 (
	   .ZN (new_n6852_),
	   .A (_net_6020) );
   NAND4_X1 g0121 (
	   .ZN (new_n6851_),
	   .A4 (new_n6850_1_),
	   .A3 (new_n6849_),
	   .A2 (new_n6847_),
	   .A1 (new_n6845_1_) );
   NAND3_X1 g0120 (
	   .ZN (new_n6850_1_),
	   .A3 (_net_6958),
	   .A2 (_net_6959),
	   .A1 (net_6934) );
   NAND3_X1 g0119 (
	   .ZN (new_n6849_),
	   .A3 (_net_6959),
	   .A2 (net_6902),
	   .A1 (new_n6848_) );
   BUF_X4 g0118 (
	   .Z (new_n6848_),
	   .A (new_n6831_1_) );
   NAND3_X1 g0117 (
	   .ZN (new_n6847_),
	   .A3 (_net_6958),
	   .A2 (net_6870),
	   .A1 (new_n6846_) );
   BUF_X4 g0116 (
	   .Z (new_n6846_),
	   .A (new_n6839_) );
   NAND2_X1 g0115 (
	   .ZN (new_n6845_1_),
	   .A2 (net_6838),
	   .A1 (new_n6844_) );
   BUF_X4 g0114 (
	   .Z (new_n6844_),
	   .A (new_n6835_) );
   AND3_X1 g0113 (
	   .ZN (new_n6843_),
	   .A3 (new_n6842_),
	   .A2 (new_n6837_),
	   .A1 (new_n6834_) );
   NAND4_X1 g0112 (
	   .ZN (new_n6842_),
	   .A4 (new_n6841_),
	   .A3 (_net_6957),
	   .A2 (net_6914),
	   .A1 (new_n6838_) );
   BUF_X4 g0111 (
	   .Z (new_n6841_),
	   .A (new_n6840_1_) );
   NOR2_X1 g0110 (
	   .ZN (new_n6840_1_),
	   .A2 (_net_6958),
	   .A1 (new_n6839_) );
   INV_X1 g0109 (
	   .ZN (new_n6839_),
	   .A (_net_6959) );
   BUF_X4 g0108 (
	   .Z (new_n6838_),
	   .A (new_n6829_) );
   NAND4_X1 g0107 (
	   .ZN (new_n6837_),
	   .A4 (new_n6836_1_),
	   .A3 (_net_6957),
	   .A2 (net_6850),
	   .A1 (new_n6830_) );
   BUF_X4 g0106 (
	   .Z (new_n6836_1_),
	   .A (new_n6835_) );
   NOR2_X1 g0105 (
	   .ZN (new_n6835_),
	   .A2 (_net_6958),
	   .A1 (_net_6959) );
   NAND4_X1 g0104 (
	   .ZN (new_n6834_),
	   .A4 (new_n6833_),
	   .A3 (net_6882),
	   .A2 (_net_6957),
	   .A1 (new_n6830_) );
   BUF_X4 g0103 (
	   .Z (new_n6833_),
	   .A (new_n6832_) );
   NOR2_X1 g0102 (
	   .ZN (new_n6832_),
	   .A2 (_net_6959),
	   .A1 (new_n6831_1_) );
   INV_X1 g0101 (
	   .ZN (new_n6831_1_),
	   .A (_net_6958) );
   BUF_X4 g0100 (
	   .Z (new_n6830_),
	   .A (new_n6829_) );
   NOR2_X1 g0099 (
	   .ZN (new_n6829_),
	   .A2 (new_n6828_),
	   .A1 (new_n6826_1_) );
   INV_X1 g0098 (
	   .ZN (new_n6828_),
	   .A (new_n6827_) );
   NOR2_X1 g0097 (
	   .ZN (new_n6827_),
	   .A2 (_net_6020),
	   .A1 (_net_6019) );
   NAND4_X1 g0096 (
	   .ZN (new_n6826_1_),
	   .A4 (_net_6017),
	   .A3 (net_6058),
	   .A2 (_net_7791),
	   .A1 (new_n6825_) );
   INV_X1 g0095 (
	   .ZN (new_n6825_),
	   .A (_net_7755) );
   MUX2_X1 g0094 (
	   .Z (n295),
	   .S (new_n6823_),
	   .B (_net_6032),
	   .A (_net_7797) );
   NAND2_X2 g0093 (
	   .ZN (new_n6823_),
	   .A2 (new_n6822_1_),
	   .A1 (new_n6820_) );
   NOR2_X1 g0092 (
	   .ZN (new_n6822_1_),
	   .A2 (x1322),
	   .A1 (new_n6821_) );
   INV_X1 g0091 (
	   .ZN (new_n6821_),
	   .A (_net_6184) );
   NOR2_X1 g0090 (
	   .ZN (new_n6820_),
	   .A2 (x1261),
	   .A1 (new_n6819_) );
   INV_X1 g0089 (
	   .ZN (new_n6819_),
	   .A (x1286) );
   CLKBUF_X1 g0088 (
	   .Z (n291),
	   .A (net_6453) );
   CLKBUF_X1 g0087 (
	   .Z (n286),
	   .A (_net_6104) );
   NAND3_X1 g0086 (
	   .ZN (n281),
	   .A3 (new_n6815_),
	   .A2 (new_n6793_1_),
	   .A1 (new_n6777_) );
   AND3_X1 g0085 (
	   .ZN (new_n6815_),
	   .A3 (new_n6814_),
	   .A2 (new_n6810_),
	   .A1 (new_n6802_) );
   NAND2_X1 g0084 (
	   .ZN (new_n6814_),
	   .A2 (_net_6082),
	   .A1 (new_n6813_1_) );
   BUF_X4 g0083 (
	   .Z (new_n6813_1_),
	   .A (new_n6812_) );
   NOR2_X1 g0082 (
	   .ZN (new_n6812_),
	   .A2 (new_n6811_),
	   .A1 (new_n6781_) );
   INV_X1 g0081 (
	   .ZN (new_n6811_),
	   .A (_net_5984) );
   NAND2_X1 g0080 (
	   .ZN (new_n6810_),
	   .A2 (new_n6809_1_),
	   .A1 (new_n6807_) );
   NOR2_X1 g0079 (
	   .ZN (new_n6809_1_),
	   .A2 (new_n6808_),
	   .A1 (new_n6760_) );
   INV_X1 g0078 (
	   .ZN (new_n6808_),
	   .A (_net_5987) );
   NAND4_X1 g0077 (
	   .ZN (new_n6807_),
	   .A4 (new_n6806_1_),
	   .A3 (new_n6805_),
	   .A2 (new_n6804_),
	   .A1 (new_n6803_) );
   NAND3_X1 g0076 (
	   .ZN (new_n6806_1_),
	   .A3 (_net_6554),
	   .A2 (net_6538),
	   .A1 (_net_6553) );
   NAND3_X1 g0075 (
	   .ZN (new_n6805_),
	   .A3 (_net_6554),
	   .A2 (net_6506),
	   .A1 (new_n6789_) );
   NAND3_X1 g0074 (
	   .ZN (new_n6804_),
	   .A3 (_net_6553),
	   .A2 (net_6474),
	   .A1 (new_n6787_) );
   NAND2_X1 g0073 (
	   .ZN (new_n6803_),
	   .A2 (net_6442),
	   .A1 (new_n6785_) );
   NAND2_X1 g0072 (
	   .ZN (new_n6802_),
	   .A2 (new_n6801_1_),
	   .A1 (new_n6798_) );
   BUF_X4 g0071 (
	   .Z (new_n6801_1_),
	   .A (new_n6800_) );
   NOR2_X1 g0070 (
	   .ZN (new_n6800_),
	   .A2 (new_n6799_),
	   .A1 (new_n6760_) );
   INV_X1 g0069 (
	   .ZN (new_n6799_),
	   .A (_net_5986) );
   NAND4_X1 g0068 (
	   .ZN (new_n6798_),
	   .A4 (new_n6797_),
	   .A3 (new_n6796_1_),
	   .A2 (new_n6795_),
	   .A1 (new_n6794_) );
   NAND3_X1 g0067 (
	   .ZN (new_n6797_),
	   .A3 (_net_6554),
	   .A2 (net_6536),
	   .A1 (_net_6553) );
   NAND3_X1 g0066 (
	   .ZN (new_n6796_1_),
	   .A3 (net_6504),
	   .A2 (_net_6554),
	   .A1 (new_n6789_) );
   NAND3_X1 g0065 (
	   .ZN (new_n6795_),
	   .A3 (net_6472),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   NAND2_X1 g0064 (
	   .ZN (new_n6794_),
	   .A2 (net_6440),
	   .A1 (new_n6785_) );
   AOI22_X1 g0063 (
	   .ZN (new_n6793_1_),
	   .B2 (new_n6792_),
	   .B1 (new_n6784_),
	   .A2 (new_n6779_1_),
	   .A1 (net_6550) );
   NAND4_X1 g0062 (
	   .ZN (new_n6792_),
	   .A4 (new_n6791_),
	   .A3 (new_n6790_),
	   .A2 (new_n6788_1_),
	   .A1 (new_n6786_) );
   NAND3_X1 g0061 (
	   .ZN (new_n6791_),
	   .A3 (net_6534),
	   .A2 (_net_6554),
	   .A1 (_net_6553) );
   NAND3_X1 g0060 (
	   .ZN (new_n6790_),
	   .A3 (_net_6554),
	   .A2 (net_6502),
	   .A1 (new_n6789_) );
   BUF_X4 g0059 (
	   .Z (new_n6789_),
	   .A (new_n6765_1_) );
   NAND3_X1 g0058 (
	   .ZN (new_n6788_1_),
	   .A3 (net_6470),
	   .A2 (_net_6553),
	   .A1 (new_n6787_) );
   BUF_X4 g0057 (
	   .Z (new_n6787_),
	   .A (new_n6773_) );
   NAND2_X1 g0056 (
	   .ZN (new_n6786_),
	   .A2 (net_6438),
	   .A1 (new_n6785_) );
   BUF_X4 g0055 (
	   .Z (new_n6785_),
	   .A (new_n6769_) );
   BUF_X4 g0054 (
	   .Z (new_n6784_),
	   .A (new_n6783_1_) );
   NOR2_X1 g0053 (
	   .ZN (new_n6783_1_),
	   .A2 (_net_6552),
	   .A1 (new_n6782_) );
   NAND3_X1 g0052 (
	   .ZN (new_n6782_),
	   .A3 (new_n6761_1_),
	   .A2 (_net_5984),
	   .A1 (new_n6781_) );
   NOR2_X1 g0051 (
	   .ZN (new_n6781_),
	   .A2 (_net_7749),
	   .A1 (new_n6780_) );
   NAND2_X1 g0050 (
	   .ZN (new_n6780_),
	   .A2 (_net_7791),
	   .A1 (net_6061) );
   NOR4_X2 g0049 (
	   .ZN (new_n6779_1_),
	   .A4 (new_n6778_),
	   .A3 (new_n6773_),
	   .A2 (new_n6762_),
	   .A1 (new_n6760_) );
   NAND2_X1 g0048 (
	   .ZN (new_n6778_),
	   .A2 (_net_6552),
	   .A1 (_net_6553) );
   AND3_X1 g0047 (
	   .ZN (new_n6777_),
	   .A3 (new_n6776_),
	   .A2 (new_n6771_),
	   .A1 (new_n6768_) );
   NAND4_X1 g0046 (
	   .ZN (new_n6776_),
	   .A4 (new_n6775_),
	   .A3 (net_6518),
	   .A2 (_net_6552),
	   .A1 (new_n6772_) );
   BUF_X4 g0045 (
	   .Z (new_n6775_),
	   .A (new_n6774_1_) );
   NOR2_X1 g0044 (
	   .ZN (new_n6774_1_),
	   .A2 (_net_6553),
	   .A1 (new_n6773_) );
   INV_X1 g0043 (
	   .ZN (new_n6773_),
	   .A (_net_6554) );
   BUF_X4 g0042 (
	   .Z (new_n6772_),
	   .A (new_n6763_) );
   NAND4_X1 g0041 (
	   .ZN (new_n6771_),
	   .A4 (new_n6770_1_),
	   .A3 (_net_6552),
	   .A2 (net_6454),
	   .A1 (new_n6764_) );
   BUF_X4 g0040 (
	   .Z (new_n6770_1_),
	   .A (new_n6769_) );
   NOR2_X1 g0039 (
	   .ZN (new_n6769_),
	   .A2 (_net_6554),
	   .A1 (_net_6553) );
   NAND4_X1 g0038 (
	   .ZN (new_n6768_),
	   .A4 (new_n6767_),
	   .A3 (_net_6552),
	   .A2 (net_6486),
	   .A1 (new_n6764_) );
   BUF_X4 g0037 (
	   .Z (new_n6767_),
	   .A (new_n6766_) );
   NOR2_X1 g0036 (
	   .ZN (new_n6766_),
	   .A2 (_net_6554),
	   .A1 (new_n6765_1_) );
   INV_X1 g0035 (
	   .ZN (new_n6765_1_),
	   .A (_net_6553) );
   BUF_X4 g0034 (
	   .Z (new_n6764_),
	   .A (new_n6763_) );
   NOR2_X1 g0033 (
	   .ZN (new_n6763_),
	   .A2 (new_n6762_),
	   .A1 (new_n6760_) );
   INV_X1 g0032 (
	   .ZN (new_n6762_),
	   .A (new_n6761_1_) );
   NOR2_X1 g0031 (
	   .ZN (new_n6761_1_),
	   .A2 (_net_5986),
	   .A1 (_net_5987) );
   NAND4_X1 g0030 (
	   .ZN (new_n6760_),
	   .A4 (_net_7791),
	   .A3 (net_6061),
	   .A2 (_net_5984),
	   .A1 (new_n6759_) );
   INV_X1 g0029 (
	   .ZN (new_n6759_),
	   .A (_net_7749) );
   CLKBUF_X1 g0028 (
	   .Z (n276),
	   .A (net_7807) );
   NAND2_X1 g0027 (
	   .ZN (n271),
	   .A2 (new_n6756_1_),
	   .A1 (new_n6754_) );
   AOI22_X1 g0026 (
	   .ZN (new_n6756_1_),
	   .B2 (_net_7576),
	   .B1 (new_n6755_),
	   .A2 (net_7608),
	   .A1 (new_n6743_) );
   BUF_X4 g0025 (
	   .Z (new_n6755_),
	   .A (new_n6750_) );
   AOI22_X1 g0024 (
	   .ZN (new_n6754_),
	   .B2 (net_7640),
	   .B1 (new_n6746_1_),
	   .A2 (new_n6749_1_),
	   .A1 (net_7672) );
   NAND2_X1 g0023 (
	   .ZN (n266),
	   .A2 (new_n6752_1_),
	   .A1 (new_n6747_) );
   AOI22_X1 g0022 (
	   .ZN (new_n6752_1_),
	   .B2 (new_n6751_),
	   .B1 (_net_7571),
	   .A2 (_net_7667),
	   .A1 (new_n6749_1_) );
   BUF_X4 g0021 (
	   .Z (new_n6751_),
	   .A (new_n6750_) );
   NOR2_X1 g0020 (
	   .ZN (new_n6750_),
	   .A2 (net_7680),
	   .A1 (_net_7681) );
   BUF_X4 g0019 (
	   .Z (new_n6749_1_),
	   .A (new_n6748_) );
   NOR2_X1 g0018 (
	   .ZN (new_n6748_),
	   .A2 (new_n6741_1_),
	   .A1 (new_n6744_) );
   AOI22_X1 g0017 (
	   .ZN (new_n6747_),
	   .B2 (_net_7635),
	   .B1 (new_n6746_1_),
	   .A2 (new_n6743_),
	   .A1 (_net_7603) );
   BUF_X4 g0016 (
	   .Z (new_n6746_1_),
	   .A (new_n6745_) );
   NOR2_X1 g0015 (
	   .ZN (new_n6745_),
	   .A2 (net_7680),
	   .A1 (new_n6744_) );
   INV_X1 g0014 (
	   .ZN (new_n6744_),
	   .A (_net_7681) );
   BUF_X4 g0013 (
	   .Z (new_n6743_),
	   .A (new_n6742_) );
   NOR2_X1 g0012 (
	   .ZN (new_n6742_),
	   .A2 (_net_7681),
	   .A1 (new_n6741_1_) );
   INV_X1 g0011 (
	   .ZN (new_n6741_1_),
	   .A (net_7680) );
   CLKBUF_X1 g0010 (
	   .Z (x77),
	   .A (_net_5851) );
   CLKBUF_X1 g0009 (
	   .Z (x114),
	   .A (_net_5856) );
   CLKBUF_X1 g0008 (
	   .Z (x101),
	   .A (_net_5854) );
   CLKBUF_X1 g0007 (
	   .Z (x106),
	   .A (_net_5855) );
   CLKBUF_X1 g0006 (
	   .Z (x96),
	   .A (_net_5853) );
   CLKBUF_X1 g0005 (
	   .Z (x63),
	   .A (_net_5850) );
   CLKBUF_X1 g0004 (
	   .Z (x145),
	   .A (x130657) );
   CLKBUF_X1 g0003 (
	   .Z (x131),
	   .A (_net_5859) );
   CLKBUF_X1 g0002 (
	   .Z (x84),
	   .A (_net_5852) );
   OR2_X1 g0001 (
	   .ZN (x30),
	   .A2 (net_6417),
	   .A1 (net_6416) );
   CLKBUF_X1 g0000 (
	   .Z (x124),
	   .A (_net_5857) );
   BUF_X4 ck_buf_22_b_0 (
	   .Z (ck_net_4_22_b_1),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_22_a_0 (
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_21_b_0 (
	   .Z (ck_net_4_21_b_1),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_21_a_0 (
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_20_b_0 (
	   .Z (ck_net_4_20_b_1),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_20_a_0 (
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_19_b_0 (
	   .Z (ck_net_4_19_b_1),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_19_a_0 (
	   .Z (ck_net_4_19_a_2),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_18_b_0 (
	   .Z (ck_net_4_18_b_1),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_18_a_0 (
	   .Z (ck_net_4_18_a_1),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_17_b_0 (
	   .Z (ck_net_4_17_b_1),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_17_a_0 (
	   .Z (ck_net_4_17_a_1),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_16_b_0 (
	   .Z (ck_net_4_16_b_1),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_16_a_0 (
	   .Z (ck_net_4_16_a_1),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_15_b_0 (
	   .Z (ck_net_4_15_b_1),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_15_a_0 (
	   .Z (ck_net_4_15_a_2),
	   .A (ck_net_1_0_b_2) );
   BUF_X4 ck_buf_14_b_0 (
	   .Z (ck_net_4_14_b_1),
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_14_a_0 (
	   .Z (ck_net_4_14_a_2),
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_13_b_0 (
	   .Z (ck_net_4_13_b_1),
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_13_a_0 (
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_12_b_0 (
	   .Z (ck_net_4_12_b_1),
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_12_a_0 (
	   .Z (ck_net_4_12_a_2),
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_11_b_0 (
	   .Z (ck_net_4_11_b_1),
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_11_a_0 (
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_10_b_0 (
	   .Z (ck_net_4_10_b_1),
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_10_a_0 (
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_9_b_0 (
	   .Z (ck_net_4_9_b_1),
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_9_a_0 (
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_8_b_0 (
	   .Z (ck_net_4_8_b_1),
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_8_a_0 (
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_7_b_0 (
	   .Z (ck_net_4_7_b_1),
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_7_a_0 (
	   .Z (ck_net_4_7_a_1),
	   .A (ck_net_1_0_a_2) );
   BUF_X4 ck_buf_0_b_0 (
	   .Z (ck_net_1_0_b_2),
	   .A (ck_net_1_0_0) );
   BUF_X4 ck_buf_0_a_0 (
	   .Z (ck_net_1_0_a_2),
	   .A (ck_net_1_0_0) );
   BUF_X4 ck_tree_0 (
	   .Z (ck_net_1_0_0),
	   .A (clk) );
endmodule

