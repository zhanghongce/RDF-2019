module ac97_ctrl (
	x977,
	x96,
	x940,
	x906,
	x889,
	x868,
	x84,
	x837,
	x821,
	x806,
	x786,
	x77,
	x765,
	x744,
	x718,
	x699,
	x681,
	x657,
	x638,
	x63,
	x620,
	x589,
	x561,
	x538,
	x522,
	x494,
	x476,
	x447,
	x420,
	x397,
	x390,
	x38,
	x379,
	x361,
	x342,
	x315,
	x30,
	x287,
	x264,
	x249,
	x234,
	x217,
	x195,
	x187,
	x1822,
	x179,
	x172,
	x1595,
	x1587,
	x1580,
	x1572,
	x1564,
	x1557,
	x1550,
	x1542,
	x1534,
	x1527,
	x1519,
	x1511,
	x1501,
	x1494,
	x149,
	x1486,
	x1479,
	x1467,
	x1459,
	x1451,
	x145,
	x1443,
	x1432,
	x1424,
	x1417,
	x1406,
	x14,
	x1398,
	x1390,
	x1382,
	x138,
	x1374,
	x1366,
	x1358,
	x1351,
	x1345,
	x1322,
	x131,
	x130657,
	x130656,
	x130655,
	x130654,
	x130653,
	x130652,
	x130651,
	x130650,
	x130649,
	x130648,
	x130647,
	x130646,
	x130645,
	x130644,
	x130643,
	x130642,
	x130641,
	x130640,
	x130639,
	x130638,
	x130637,
	x130636,
	x130635,
	x130634,
	x130633,
	x130632,
	x130631,
	x130630,
	x130629,
	x1286,
	x1261,
	x124,
	x1231,
	x1215,
	x1209,
	x1203,
	x1193,
	x1155,
	x114,
	x1126,
	x1101,
	x1062,
	x106,
	x1034,
	x101,
	x1006,
	x0,
	clk);
   input x977;
   output x96;
   input x940;
   input x906;
   input x889;
   input x868;
   output x84;
   input x837;
   input x821;
   input x806;
   output x786;
   output x77;
   output x765;
   output x744;
   output x718;
   output x699;
   output x681;
   output x657;
   output x638;
   output x63;
   output x620;
   output x589;
   output x561;
   output x538;
   output x522;
   output x494;
   output x476;
   output x447;
   output x420;
   output x397;
   output x390;
   output x38;
   output x379;
   output x361;
   output x342;
   output x315;
   output x30;
   output x287;
   output x264;
   output x249;
   output x234;
   output x217;
   output x195;
   output x187;
   input x1822;
   output x179;
   output x172;
   input x1595;
   input x1587;
   input x1580;
   input x1572;
   input x1564;
   input x1557;
   input x1550;
   input x1542;
   input x1534;
   input x1527;
   input x1519;
   input x1511;
   input x1501;
   input x1494;
   output x149;
   input x1486;
   input x1479;
   input x1467;
   input x1459;
   input x1451;
   output x145;
   input x1443;
   input x1432;
   input x1424;
   input x1417;
   input x1406;
   output x14;
   input x1398;
   input x1390;
   input x1382;
   output x138;
   input x1374;
   input x1366;
   input x1358;
   input x1351;
   input x1345;
   input x1322;
   output x131;
   input x130657;
   input x130656;
   input x130655;
   input x130654;
   input x130653;
   input x130652;
   input x130651;
   input x130650;
   input x130649;
   input x130648;
   input x130647;
   input x130646;
   input x130645;
   input x130644;
   input x130643;
   input x130642;
   input x130641;
   input x130640;
   input x130639;
   input x130638;
   input x130637;
   input x130636;
   input x130635;
   input x130634;
   input x130633;
   input x130632;
   input x130631;
   input x130630;
   input x130629;
   input x1286;
   input x1261;
   output x124;
   input x1231;
   input x1215;
   input x1209;
   input x1203;
   input x1193;
   input x1155;
   output x114;
   input x1126;
   input x1101;
   input x1062;
   output x106;
   input x1034;
   output x101;
   input x1006;
   output x0;
   input clk;

   // Internal wires
   wire x977;
   wire x96;
   wire x940;
   wire x906;
   wire x889;
   wire x868;
   wire x84;
   wire x837;
   wire x821;
   wire x806;
   wire x786;
   wire x77;
   wire x765;
   wire x744;
   wire x718;
   wire x699;
   wire x681;
   wire x657;
   wire x638;
   wire x63;
   wire x620;
   wire x589;
   wire x561;
   wire x538;
   wire x522;
   wire x494;
   wire x476;
   wire x447;
   wire x420;
   wire x397;
   wire x390;
   wire x38;
   wire x379;
   wire x361;
   wire x342;
   wire x315;
   wire x30;
   wire x287;
   wire x264;
   wire x249;
   wire x234;
   wire x217;
   wire x195;
   wire x187;
   wire x1822;
   wire x179;
   wire x172;
   wire x1595;
   wire x1587;
   wire x1580;
   wire x1572;
   wire x1564;
   wire x1557;
   wire x1550;
   wire x1542;
   wire x1534;
   wire x1527;
   wire x1519;
   wire x1511;
   wire x1501;
   wire x1494;
   wire x149;
   wire x1486;
   wire x1479;
   wire x1467;
   wire x1459;
   wire x1451;
   wire x145;
   wire x1443;
   wire x1432;
   wire x1424;
   wire x1417;
   wire x1406;
   wire x14;
   wire x1398;
   wire x1390;
   wire x1382;
   wire x138;
   wire x1374;
   wire x1366;
   wire x1358;
   wire x1351;
   wire x1345;
   wire x1322;
   wire x131;
   wire x130657;
   wire x130656;
   wire x130655;
   wire x130654;
   wire x130653;
   wire x130652;
   wire x130651;
   wire x130650;
   wire x130649;
   wire x130648;
   wire x130647;
   wire x130646;
   wire x130645;
   wire x130644;
   wire x130643;
   wire x130642;
   wire x130641;
   wire x130640;
   wire x130639;
   wire x130638;
   wire x130637;
   wire x130636;
   wire x130635;
   wire x130634;
   wire x130633;
   wire x130632;
   wire x130631;
   wire x130630;
   wire x130629;
   wire x1286;
   wire x1261;
   wire x124;
   wire x1231;
   wire x1215;
   wire x1209;
   wire x1203;
   wire x1193;
   wire x1155;
   wire x114;
   wire x1126;
   wire x1101;
   wire x1062;
   wire x106;
   wire x1034;
   wire x101;
   wire x1006;
   wire x0;
   wire new_n9999_;
   wire new_n9998_;
   wire new_n9997_1_;
   wire new_n9996_;
   wire new_n9995_;
   wire new_n9994_;
   wire new_n9993_;
   wire new_n9992_1_;
   wire new_n9991_;
   wire new_n9990_;
   wire new_n9989_;
   wire new_n9988_1_;
   wire new_n9987_;
   wire new_n9986_;
   wire new_n9985_1_;
   wire new_n9984_;
   wire new_n9983_;
   wire new_n9982_;
   wire new_n9981_1_;
   wire new_n9976_1_;
   wire new_n9975_;
   wire new_n9974_;
   wire new_n9973_;
   wire new_n9972_;
   wire new_n9971_1_;
   wire new_n9970_;
   wire new_n9969_;
   wire new_n9968_;
   wire new_n9967_;
   wire new_n9966_1_;
   wire new_n9965_;
   wire new_n9964_;
   wire new_n9963_;
   wire new_n9951_;
   wire new_n9950_;
   wire new_n9949_1_;
   wire new_n9939_1_;
   wire new_n9938_;
   wire new_n9935_1_;
   wire new_n9934_;
   wire new_n9933_;
   wire new_n9928_;
   wire new_n9927_;
   wire new_n9920_;
   wire new_n9919_;
   wire new_n9918_1_;
   wire new_n9917_;
   wire new_n9916_;
   wire new_n9915_;
   wire new_n9914_1_;
   wire new_n9910_;
   wire new_n9909_;
   wire new_n9908_;
   wire new_n9903_;
   wire new_n9902_1_;
   wire new_n9901_;
   wire new_n9900_;
   wire new_n9885_1_;
   wire new_n9883_;
   wire new_n9881_;
   wire new_n9876_;
   wire new_n9875_1_;
   wire new_n9874_;
   wire new_n9873_;
   wire new_n9872_;
   wire new_n9871_1_;
   wire new_n9870_;
   wire new_n9869_;
   wire new_n9868_;
   wire new_n9867_1_;
   wire new_n9866_;
   wire new_n9865_;
   wire new_n9857_;
   wire new_n9856_;
   wire new_n9855_;
   wire new_n9854_;
   wire new_n9853_1_;
   wire new_n9852_;
   wire new_n9851_;
   wire new_n9850_;
   wire new_n9849_1_;
   wire new_n9848_;
   wire new_n9847_;
   wire new_n9846_;
   wire new_n9844_1_;
   wire new_n9839_;
   wire new_n9838_;
   wire new_n9835_;
   wire new_n9834_;
   wire new_n9832_;
   wire new_n9831_;
   wire new_n9830_;
   wire new_n9829_;
   wire new_n9828_1_;
   wire new_n9826_;
   wire new_n9825_;
   wire new_n9822_;
   wire new_n9821_;
   wire new_n9813_;
   wire new_n9812_;
   wire new_n9810_;
   wire new_n9805_1_;
   wire new_n9804_;
   wire new_n9803_;
   wire new_n9798_;
   wire new_n9797_;
   wire new_n9794_;
   wire new_n9793_;
   wire new_n9791_;
   wire new_n9790_;
   wire new_n9789_;
   wire new_n9788_;
   wire new_n9787_1_;
   wire new_n9786_;
   wire new_n9785_;
   wire new_n9784_;
   wire new_n9783_1_;
   wire new_n9782_;
   wire new_n9781_;
   wire new_n9780_;
   wire new_n9779_;
   wire new_n9778_1_;
   wire new_n9777_;
   wire new_n9776_;
   wire new_n9775_;
   wire new_n9774_;
   wire new_n9773_1_;
   wire new_n9768_1_;
   wire new_n9767_;
   wire new_n9765_;
   wire new_n9764_;
   wire new_n9763_1_;
   wire new_n9762_;
   wire new_n9761_;
   wire new_n9760_;
   wire new_n9759_;
   wire new_n9758_1_;
   wire new_n9757_;
   wire new_n9755_;
   wire new_n9752_;
   wire new_n9747_;
   wire new_n9746_1_;
   wire new_n9745_;
   wire new_n9744_;
   wire new_n9743_;
   wire new_n9742_1_;
   wire new_n9741_;
   wire new_n9736_;
   wire new_n9735_;
   wire new_n9732_;
   wire new_n9731_;
   wire new_n9730_;
   wire new_n9729_1_;
   wire new_n9724_1_;
   wire new_n9723_;
   wire new_n9722_;
   wire new_n9721_;
   wire new_n9720_;
   wire new_n9718_;
   wire new_n9717_;
   wire new_n9708_;
   wire new_n9707_;
   wire new_n9703_;
   wire new_n9702_;
   wire new_n9694_;
   wire new_n9693_;
   wire new_n9686_;
   wire new_n9685_;
   wire new_n9684_;
   wire new_n9683_1_;
   wire new_n9682_;
   wire new_n9679_;
   wire new_n9678_1_;
   wire new_n9677_;
   wire new_n9676_;
   wire new_n9675_;
   wire new_n9674_;
   wire new_n9673_1_;
   wire new_n9670_;
   wire new_n9669_;
   wire new_n9668_1_;
   wire new_n9667_;
   wire new_n9666_;
   wire new_n9665_;
   wire new_n9664_1_;
   wire new_n9662_;
   wire new_n9661_;
   wire new_n9659_;
   wire new_n9651_1_;
   wire new_n9650_;
   wire new_n9649_;
   wire new_n9648_;
   wire new_n9647_1_;
   wire new_n9646_;
   wire new_n9645_;
   wire new_n9644_;
   wire new_n9643_;
   wire new_n9637_;
   wire new_n9636_;
   wire new_n9635_;
   wire new_n9634_;
   wire new_n9633_1_;
   wire new_n9632_;
   wire new_n9631_;
   wire new_n9630_;
   wire new_n9629_;
   wire new_n9628_1_;
   wire new_n9627_;
   wire new_n9623_;
   wire new_n9620_1_;
   wire new_n9619_;
   wire new_n9618_;
   wire new_n9613_;
   wire new_n9612_;
   wire new_n9611_1_;
   wire new_n9610_;
   wire new_n9608_;
   wire new_n9607_;
   wire new_n9604_;
   wire new_n9602_1_;
   wire new_n9601_;
   wire new_n9594_;
   wire new_n9593_;
   wire new_n9591_;
   wire new_n9590_;
   wire new_n9587_;
   wire new_n9586_;
   wire new_n9584_;
   wire new_n9583_1_;
   wire new_n9581_;
   wire new_n9580_;
   wire new_n9574_1_;
   wire new_n9573_;
   wire new_n9571_;
   wire new_n9570_;
   wire new_n9569_1_;
   wire new_n9562_;
   wire new_n9561_;
   wire new_n9560_;
   wire new_n9559_1_;
   wire new_n9558_;
   wire new_n9546_1_;
   wire new_n9541_1_;
   wire new_n9540_;
   wire new_n9539_;
   wire new_n9538_;
   wire new_n9537_1_;
   wire new_n9536_;
   wire new_n9531_;
   wire new_n9530_;
   wire new_n9529_;
   wire new_n9528_1_;
   wire new_n9527_;
   wire new_n9526_;
   wire new_n9525_1_;
   wire new_n9524_;
   wire new_n9523_;
   wire new_n9522_;
   wire new_n9520_1_;
   wire new_n9517_1_;
   wire new_n9516_;
   wire new_n9509_;
   wire new_n9508_;
   wire new_n9507_1_;
   wire new_n9504_;
   wire new_n9503_;
   wire new_n9502_1_;
   wire new_n9501_;
   wire new_n9498_;
   wire new_n9497_1_;
   wire new_n9496_;
   wire new_n9495_;
   wire new_n9494_;
   wire new_n9493_;
   wire new_n9492_1_;
   wire new_n9491_;
   wire new_n9490_;
   wire new_n9489_;
   wire new_n9488_;
   wire new_n9487_1_;
   wire new_n9486_;
   wire new_n9485_;
   wire new_n9484_;
   wire new_n9481_;
   wire new_n9480_;
   wire new_n9478_1_;
   wire new_n9477_;
   wire new_n9469_;
   wire new_n9468_;
   wire new_n9467_1_;
   wire new_n9465_;
   wire new_n9464_;
   wire new_n9463_;
   wire new_n9462_1_;
   wire new_n9458_;
   wire new_n9457_;
   wire new_n9453_;
   wire new_n9452_;
   wire new_n9451_;
   wire new_n9450_;
   wire new_n9449_1_;
   wire new_n9448_;
   wire new_n9447_;
   wire new_n9446_;
   wire new_n9445_1_;
   wire new_n9442_;
   wire new_n9441_1_;
   wire new_n9440_;
   wire new_n9439_;
   wire new_n9438_;
   wire new_n9436_1_;
   wire new_n9435_;
   wire new_n9434_;
   wire new_n9433_;
   wire new_n9428_1_;
   wire new_n9427_;
   wire new_n9426_;
   wire new_n9421_;
   wire new_n9420_1_;
   wire new_n9417_;
   wire new_n9416_;
   wire new_n9405_1_;
   wire new_n9404_;
   wire new_n9403_;
   wire new_n9401_;
   wire new_n9400_;
   wire new_n9393_1_;
   wire new_n9392_;
   wire new_n9391_;
   wire new_n9387_;
   wire new_n9385_1_;
   wire new_n9384_;
   wire new_n9381_1_;
   wire new_n9380_;
   wire new_n9378_;
   wire new_n9377_1_;
   wire new_n9376_;
   wire new_n9375_;
   wire new_n9374_;
   wire new_n9371_;
   wire new_n9370_1_;
   wire new_n9367_;
   wire new_n9366_;
   wire new_n9360_;
   wire new_n9359_;
   wire new_n9358_;
   wire new_n9357_;
   wire new_n9356_1_;
   wire new_n9355_;
   wire new_n9354_;
   wire new_n9351_;
   wire new_n9349_;
   wire new_n9348_1_;
   wire new_n9347_;
   wire new_n9345_;
   wire new_n9344_;
   wire new_n9343_1_;
   wire new_n9342_;
   wire new_n9341_;
   wire new_n9340_;
   wire new_n9339_1_;
   wire new_n9338_;
   wire new_n9333_;
   wire new_n9332_;
   wire new_n9331_;
   wire new_n9330_1_;
   wire new_n9329_;
   wire new_n9328_;
   wire new_n9327_;
   wire new_n9326_1_;
   wire new_n9325_;
   wire new_n9324_;
   wire new_n9323_;
   wire new_n9322_;
   wire new_n9321_1_;
   wire new_n9320_;
   wire new_n9316_1_;
   wire new_n9315_;
   wire new_n9311_;
   wire new_n9310_;
   wire new_n9308_;
   wire new_n9307_1_;
   wire new_n9306_;
   wire new_n9305_;
   wire new_n9304_;
   wire new_n9303_;
   wire new_n9289_;
   wire new_n9288_;
   wire new_n9285_;
   wire new_n9284_;
   wire new_n9283_;
   wire new_n9282_1_;
   wire new_n9281_;
   wire new_n9280_;
   wire new_n9279_;
   wire new_n9278_;
   wire new_n9277_1_;
   wire new_n9276_;
   wire new_n9275_;
   wire new_n9274_;
   wire new_n9273_;
   wire new_n9272_1_;
   wire new_n9271_;
   wire new_n9270_;
   wire new_n9269_;
   wire new_n9268_;
   wire new_n9267_1_;
   wire new_n9262_;
   wire new_n9261_;
   wire new_n9257_;
   wire new_n9256_;
   wire new_n9255_;
   wire new_n9254_1_;
   wire new_n9253_;
   wire new_n9252_;
   wire new_n9251_;
   wire new_n9250_1_;
   wire new_n9249_;
   wire new_n9248_;
   wire new_n9247_;
   wire new_n9243_;
   wire new_n9242_1_;
   wire new_n9241_;
   wire new_n9240_;
   wire new_n9239_;
   wire new_n9238_1_;
   wire new_n9237_;
   wire new_n9236_;
   wire new_n9235_;
   wire new_n9234_;
   wire new_n9233_1_;
   wire new_n9232_;
   wire new_n9231_;
   wire new_n9230_;
   wire new_n9228_1_;
   wire new_n9227_;
   wire new_n9226_;
   wire new_n9225_1_;
   wire new_n9224_;
   wire new_n9223_;
   wire new_n9222_;
   wire new_n9221_;
   wire new_n9220_1_;
   wire new_n9219_;
   wire new_n9218_;
   wire new_n9217_;
   wire new_n9216_;
   wire new_n9215_1_;
   wire new_n9211_1_;
   wire new_n9210_;
   wire new_n9205_;
   wire new_n9204_;
   wire new_n9203_;
   wire new_n9197_;
   wire new_n9196_1_;
   wire new_n9195_;
   wire new_n9193_;
   wire new_n9192_1_;
   wire new_n9191_;
   wire new_n9190_;
   wire new_n9189_;
   wire new_n9188_;
   wire new_n9187_1_;
   wire new_n9186_;
   wire new_n9185_;
   wire new_n9184_;
   wire new_n9183_;
   wire new_n9182_1_;
   wire new_n9181_;
   wire new_n9180_;
   wire new_n9179_;
   wire new_n9178_1_;
   wire new_n9177_;
   wire new_n9176_;
   wire new_n9175_;
   wire new_n9174_;
   wire new_n9173_1_;
   wire new_n9172_;
   wire new_n9171_;
   wire new_n9170_;
   wire new_n9163_;
   wire new_n9162_;
   wire new_n9161_;
   wire new_n9160_1_;
   wire new_n9159_;
   wire new_n9158_;
   wire new_n9156_1_;
   wire new_n9155_;
   wire new_n9149_;
   wire new_n9148_;
   wire new_n9147_;
   wire new_n9146_1_;
   wire new_n9145_;
   wire new_n9144_;
   wire new_n9143_1_;
   wire new_n9142_;
   wire new_n9141_;
   wire new_n9140_;
   wire new_n9139_;
   wire new_n9138_1_;
   wire new_n9137_;
   wire new_n9136_;
   wire new_n9135_;
   wire new_n9127_;
   wire new_n9126_;
   wire new_n9125_;
   wire new_n9124_1_;
   wire new_n9123_;
   wire new_n9122_;
   wire new_n9121_;
   wire new_n9120_1_;
   wire new_n9119_;
   wire new_n9118_;
   wire new_n9117_;
   wire new_n9116_;
   wire new_n9113_;
   wire new_n9112_;
   wire new_n9111_;
   wire new_n9110_1_;
   wire new_n9109_;
   wire new_n9108_;
   wire new_n9107_;
   wire new_n9106_1_;
   wire new_n9105_;
   wire new_n9103_;
   wire new_n9102_;
   wire new_n9098_;
   wire new_n9097_;
   wire new_n9096_1_;
   wire new_n9095_;
   wire new_n9094_;
   wire new_n9093_;
   wire new_n9092_;
   wire new_n9091_1_;
   wire new_n9090_;
   wire new_n9089_;
   wire new_n9088_;
   wire new_n9087_;
   wire new_n9086_1_;
   wire new_n9085_;
   wire new_n9084_;
   wire new_n9083_;
   wire new_n9082_1_;
   wire new_n9081_;
   wire new_n9080_;
   wire new_n9073_;
   wire new_n9072_;
   wire new_n9071_;
   wire new_n9070_;
   wire new_n9069_1_;
   wire new_n9068_;
   wire new_n9067_;
   wire new_n9066_;
   wire new_n9065_1_;
   wire new_n9058_;
   wire new_n9057_1_;
   wire new_n9056_;
   wire new_n9055_;
   wire new_n9054_;
   wire new_n9053_;
   wire new_n9052_1_;
   wire new_n9051_;
   wire new_n9050_;
   wire new_n9049_;
   wire new_n9048_;
   wire new_n9047_1_;
   wire new_n9046_;
   wire new_n9045_;
   wire new_n9042_1_;
   wire new_n9039_;
   wire new_n9038_;
   wire new_n9037_1_;
   wire new_n9036_;
   wire new_n9035_;
   wire new_n9033_;
   wire new_n9032_;
   wire new_n9031_;
   wire new_n9030_1_;
   wire new_n9029_;
   wire new_n9028_;
   wire new_n9027_;
   wire new_n9026_;
   wire new_n9025_1_;
   wire new_n9024_;
   wire new_n9023_;
   wire new_n9022_1_;
   wire new_n9021_;
   wire new_n9020_;
   wire new_n9018_;
   wire new_n9017_1_;
   wire new_n9014_1_;
   wire new_n9013_;
   wire new_n9012_;
   wire new_n9009_;
   wire new_n9008_;
   wire new_n9003_;
   wire new_n9002_;
   wire new_n9001_;
   wire new_n8997_;
   wire new_n8996_;
   wire new_n8991_;
   wire new_n8990_1_;
   wire new_n8985_;
   wire new_n8984_;
   wire new_n8973_;
   wire new_n8972_;
   wire new_n8969_;
   wire new_n8968_;
   wire new_n8964_;
   wire new_n8963_1_;
   wire new_n8962_;
   wire new_n8959_;
   wire new_n8958_1_;
   wire new_n8957_;
   wire new_n8948_1_;
   wire new_n8947_;
   wire new_n8945_;
   wire new_n8944_;
   wire new_n8940_;
   wire new_n8939_1_;
   wire new_n8938_;
   wire new_n8937_;
   wire new_n8936_;
   wire new_n8935_;
   wire new_n8934_1_;
   wire new_n8933_;
   wire new_n8932_;
   wire new_n8931_1_;
   wire new_n8930_;
   wire new_n8929_;
   wire new_n8928_;
   wire new_n8927_;
   wire new_n8925_;
   wire new_n8924_;
   wire new_n8923_;
   wire new_n8922_1_;
   wire new_n8921_;
   wire new_n8920_;
   wire new_n8919_;
   wire new_n8916_;
   wire new_n8915_;
   wire new_n8913_;
   wire new_n8912_1_;
   wire new_n8911_;
   wire new_n8909_;
   wire new_n8908_1_;
   wire new_n8907_;
   wire new_n8905_;
   wire new_n8899_1_;
   wire new_n8898_;
   wire new_n8897_;
   wire new_n8888_;
   wire new_n8887_;
   wire new_n8886_1_;
   wire new_n8885_;
   wire new_n8884_;
   wire new_n8883_;
   wire new_n8882_1_;
   wire new_n8881_;
   wire new_n8880_;
   wire new_n8879_;
   wire new_n8878_;
   wire new_n8873_1_;
   wire new_n8872_;
   wire new_n8861_;
   wire new_n8860_1_;
   wire new_n8859_;
   wire new_n8858_;
   wire new_n8857_;
   wire new_n8854_;
   wire new_n8853_;
   wire new_n8852_;
   wire new_n8851_;
   wire new_n8848_;
   wire new_n8846_;
   wire new_n8845_1_;
   wire new_n8844_;
   wire new_n8843_;
   wire new_n8842_;
   wire new_n8841_;
   wire new_n8840_1_;
   wire new_n8839_;
   wire new_n8838_;
   wire new_n8837_;
   wire new_n8836_;
   wire new_n8835_1_;
   wire new_n8834_;
   wire new_n8833_;
   wire new_n8832_;
   wire new_n8831_1_;
   wire new_n8830_;
   wire new_n8829_;
   wire new_n8828_;
   wire new_n8822_;
   wire new_n8821_;
   wire new_n8817_;
   wire new_n8816_;
   wire new_n8810_;
   wire new_n8805_1_;
   wire new_n8804_;
   wire new_n8803_;
   wire new_n8802_;
   wire new_n8801_;
   wire new_n8800_1_;
   wire new_n8799_;
   wire new_n8798_;
   wire new_n8797_1_;
   wire new_n8796_;
   wire new_n8795_;
   wire new_n8794_;
   wire new_n8793_1_;
   wire new_n8792_;
   wire new_n8790_;
   wire new_n8789_;
   wire new_n8788_1_;
   wire new_n8782_;
   wire new_n8781_;
   wire new_n8780_1_;
   wire new_n8779_;
   wire new_n8778_;
   wire new_n8774_;
   wire new_n8773_;
   wire new_n8767_1_;
   wire new_n8766_;
   wire new_n8765_;
   wire new_n8764_;
   wire new_n8761_;
   wire new_n8760_;
   wire new_n8759_;
   wire new_n8758_;
   wire new_n8757_1_;
   wire new_n8756_;
   wire new_n8755_;
   wire new_n8754_;
   wire new_n8753_1_;
   wire new_n8747_;
   wire new_n8746_;
   wire new_n8745_;
   wire new_n8744_;
   wire new_n8743_1_;
   wire new_n8742_;
   wire new_n8741_;
   wire new_n8740_;
   wire new_n8739_1_;
   wire new_n8738_;
   wire new_n8737_;
   wire new_n8736_;
   wire new_n8735_;
   wire new_n8734_1_;
   wire new_n8733_;
   wire new_n8732_;
   wire new_n8731_;
   wire new_n8730_1_;
   wire new_n8729_;
   wire new_n8728_;
   wire new_n8727_;
   wire new_n8726_;
   wire new_n8725_1_;
   wire new_n8724_;
   wire new_n8723_;
   wire new_n8719_;
   wire new_n8718_;
   wire new_n8717_;
   wire new_n8713_;
   wire new_n8712_;
   wire new_n8700_;
   wire new_n8698_1_;
   wire new_n8696_;
   wire new_n8695_;
   wire new_n8694_1_;
   wire new_n8692_;
   wire new_n8691_;
   wire new_n8690_;
   wire new_n8687_;
   wire new_n8686_;
   wire new_n8685_1_;
   wire new_n8681_1_;
   wire new_n8680_;
   wire new_n8679_;
   wire new_n8678_;
   wire new_n8677_;
   wire new_n8675_;
   wire new_n8671_1_;
   wire new_n8670_;
   wire new_n8669_;
   wire new_n8668_;
   wire new_n8667_;
   wire new_n8666_1_;
   wire new_n8665_;
   wire new_n8664_;
   wire new_n8663_;
   wire new_n8662_1_;
   wire new_n8661_;
   wire new_n8660_;
   wire new_n8659_;
   wire new_n8658_1_;
   wire new_n8657_;
   wire new_n8656_;
   wire new_n8655_;
   wire new_n8654_1_;
   wire new_n8653_;
   wire new_n8652_;
   wire new_n8651_;
   wire new_n8650_1_;
   wire new_n8649_;
   wire new_n8648_;
   wire new_n8646_;
   wire new_n8645_1_;
   wire new_n8643_;
   wire new_n8642_;
   wire new_n8641_1_;
   wire new_n8637_1_;
   wire new_n8636_;
   wire new_n8629_;
   wire new_n8628_1_;
   wire new_n8626_;
   wire new_n8625_1_;
   wire new_n8622_;
   wire new_n8621_1_;
   wire new_n8620_;
   wire new_n8619_;
   wire new_n8618_;
   wire new_n8617_;
   wire new_n8616_1_;
   wire new_n8615_;
   wire new_n8614_;
   wire new_n8613_;
   wire new_n8612_1_;
   wire new_n8611_;
   wire new_n8610_;
   wire new_n8609_;
   wire new_n8608_;
   wire new_n8601_;
   wire new_n8600_;
   wire new_n8599_;
   wire new_n8598_1_;
   wire new_n8597_;
   wire new_n8596_;
   wire new_n8594_;
   wire new_n8593_1_;
   wire new_n8592_;
   wire new_n8591_;
   wire new_n8587_;
   wire new_n8586_;
   wire new_n8581_;
   wire new_n8580_;
   wire new_n8579_;
   wire new_n8578_1_;
   wire new_n8577_;
   wire new_n8576_;
   wire new_n8575_1_;
   wire new_n8574_;
   wire new_n8573_;
   wire new_n8572_;
   wire new_n8571_;
   wire new_n8570_1_;
   wire new_n8569_;
   wire new_n8568_;
   wire new_n8566_;
   wire new_n8565_1_;
   wire new_n8561_1_;
   wire new_n8560_;
   wire new_n8559_;
   wire new_n8556_;
   wire new_n8555_;
   wire new_n8554_;
   wire new_n8553_;
   wire new_n8552_1_;
   wire new_n8551_;
   wire new_n8550_;
   wire new_n8549_1_;
   wire new_n8548_;
   wire new_n8547_;
   wire new_n8546_;
   wire new_n8545_;
   wire new_n8543_;
   wire new_n8541_;
   wire new_n8540_1_;
   wire new_n8536_;
   wire new_n8535_1_;
   wire new_n8534_;
   wire new_n8533_;
   wire new_n8532_;
   wire new_n8531_1_;
   wire new_n8530_;
   wire new_n8529_;
   wire new_n8528_;
   wire new_n8527_;
   wire new_n8526_1_;
   wire new_n8525_;
   wire new_n8524_;
   wire new_n8523_;
   wire new_n8522_1_;
   wire new_n8521_;
   wire new_n8520_;
   wire new_n8519_;
   wire new_n8518_;
   wire new_n8517_1_;
   wire new_n8516_;
   wire new_n8515_;
   wire new_n8514_;
   wire new_n8513_1_;
   wire new_n8505_;
   wire new_n8503_;
   wire new_n8502_;
   wire new_n8501_;
   wire new_n8500_;
   wire new_n8499_1_;
   wire new_n8498_;
   wire new_n8497_;
   wire new_n8496_;
   wire new_n8495_;
   wire new_n8494_1_;
   wire new_n8493_;
   wire new_n8492_;
   wire new_n8491_1_;
   wire new_n8490_;
   wire new_n8489_;
   wire new_n8488_;
   wire new_n8487_;
   wire new_n8486_1_;
   wire new_n8485_;
   wire new_n8484_;
   wire new_n8483_;
   wire new_n8482_;
   wire new_n8481_1_;
   wire new_n8480_;
   wire new_n8475_;
   wire new_n8474_;
   wire new_n8473_;
   wire new_n8469_;
   wire new_n8468_;
   wire new_n8463_;
   wire new_n8461_;
   wire new_n8460_;
   wire new_n8459_1_;
   wire new_n8458_;
   wire new_n8457_;
   wire new_n8456_;
   wire new_n8455_1_;
   wire new_n8454_;
   wire new_n8453_;
   wire new_n8452_;
   wire new_n8451_1_;
   wire new_n8450_;
   wire new_n8449_;
   wire new_n8448_;
   wire new_n8447_1_;
   wire new_n8446_;
   wire new_n8445_;
   wire new_n8444_;
   wire new_n8443_1_;
   wire new_n8441_;
   wire new_n8440_;
   wire new_n8439_;
   wire new_n8438_1_;
   wire new_n8436_;
   wire new_n8435_1_;
   wire new_n8431_;
   wire new_n8430_1_;
   wire new_n8429_;
   wire new_n8428_;
   wire new_n8427_;
   wire new_n8426_1_;
   wire new_n8425_;
   wire new_n8424_;
   wire new_n8423_;
   wire new_n8422_1_;
   wire new_n8421_;
   wire new_n8420_;
   wire new_n8419_;
   wire new_n8418_1_;
   wire new_n8416_;
   wire new_n8415_1_;
   wire new_n8412_;
   wire new_n8411_;
   wire new_n8410_1_;
   wire new_n8407_;
   wire new_n8406_;
   wire new_n8405_1_;
   wire new_n8404_;
   wire new_n8403_;
   wire new_n8402_;
   wire new_n8401_1_;
   wire new_n8400_;
   wire new_n8396_1_;
   wire new_n8395_;
   wire new_n8394_;
   wire new_n8393_;
   wire new_n8392_1_;
   wire new_n8391_;
   wire new_n8390_;
   wire new_n8389_;
   wire new_n8387_1_;
   wire new_n8386_;
   wire new_n8383_;
   wire new_n8382_1_;
   wire new_n8381_;
   wire new_n8380_;
   wire new_n8379_;
   wire new_n8377_1_;
   wire new_n8376_;
   wire new_n8375_;
   wire new_n8374_;
   wire new_n8373_;
   wire new_n8372_1_;
   wire new_n8371_;
   wire new_n8370_;
   wire new_n8369_;
   wire new_n8368_;
   wire new_n8367_1_;
   wire new_n8366_;
   wire new_n8365_;
   wire new_n8364_;
   wire new_n8363_;
   wire new_n8362_1_;
   wire new_n8361_;
   wire new_n8360_;
   wire new_n8359_1_;
   wire new_n8358_;
   wire new_n8357_;
   wire new_n8356_;
   wire new_n8355_;
   wire new_n8354_1_;
   wire new_n8350_1_;
   wire new_n8349_;
   wire new_n8348_;
   wire new_n8347_;
   wire new_n8346_;
   wire new_n8345_1_;
   wire new_n8344_;
   wire new_n8343_;
   wire new_n8342_;
   wire new_n8341_;
   wire new_n8339_;
   wire new_n8338_;
   wire new_n8336_;
   wire new_n8335_;
   wire new_n8334_1_;
   wire new_n8327_;
   wire new_n8326_;
   wire new_n8325_;
   wire new_n8324_1_;
   wire new_n8307_1_;
   wire new_n8306_;
   wire new_n8305_;
   wire new_n8304_;
   wire new_n8303_1_;
   wire new_n8301_;
   wire new_n8300_;
   wire new_n8299_1_;
   wire new_n8298_;
   wire new_n8297_;
   wire new_n8296_;
   wire new_n8294_1_;
   wire new_n8293_;
   wire new_n8292_;
   wire new_n8291_;
   wire new_n8289_1_;
   wire new_n8288_;
   wire new_n8285_;
   wire new_n8284_1_;
   wire new_n8282_;
   wire new_n8281_;
   wire new_n8280_1_;
   wire new_n8276_1_;
   wire new_n8275_;
   wire new_n8274_;
   wire new_n8273_;
   wire new_n8272_;
   wire new_n8271_1_;
   wire new_n8270_;
   wire new_n8269_;
   wire new_n8267_;
   wire new_n8266_1_;
   wire new_n8265_;
   wire new_n8263_;
   wire new_n8262_1_;
   wire new_n8254_;
   wire new_n8253_1_;
   wire new_n8252_;
   wire new_n8251_;
   wire new_n8250_;
   wire new_n8249_1_;
   wire new_n8248_;
   wire new_n8247_;
   wire new_n8246_;
   wire new_n8245_1_;
   wire new_n8244_;
   wire new_n8243_;
   wire new_n8234_;
   wire new_n8233_;
   wire new_n8231_;
   wire new_n8230_;
   wire new_n8229_;
   wire new_n8228_1_;
   wire new_n8225_;
   wire new_n8224_1_;
   wire new_n8221_;
   wire new_n8220_1_;
   wire new_n8219_;
   wire new_n8218_;
   wire new_n8217_;
   wire new_n8216_1_;
   wire new_n8215_;
   wire new_n8214_;
   wire new_n8212_;
   wire new_n8211_1_;
   wire new_n8210_;
   wire new_n8209_;
   wire new_n8208_;
   wire new_n8207_;
   wire new_n8206_1_;
   wire new_n8205_;
   wire new_n8204_;
   wire new_n8203_;
   wire new_n8202_1_;
   wire new_n8201_;
   wire new_n8200_;
   wire new_n8199_;
   wire new_n8198_;
   wire new_n8197_1_;
   wire new_n8193_;
   wire new_n8192_1_;
   wire new_n8191_;
   wire new_n8188_1_;
   wire new_n8187_;
   wire new_n8186_;
   wire new_n8185_;
   wire new_n8184_;
   wire new_n8183_1_;
   wire new_n8181_;
   wire new_n8180_;
   wire new_n8179_1_;
   wire new_n8178_;
   wire new_n8177_;
   wire new_n8176_;
   wire new_n8175_;
   wire new_n8174_1_;
   wire new_n8173_;
   wire new_n8172_;
   wire new_n8171_;
   wire new_n8170_1_;
   wire new_n8169_;
   wire new_n8168_;
   wire new_n8167_;
   wire new_n8166_1_;
   wire new_n8165_;
   wire new_n8164_;
   wire new_n8163_;
   wire new_n8162_;
   wire new_n8161_1_;
   wire new_n8160_;
   wire new_n8159_;
   wire new_n8158_;
   wire new_n8157_;
   wire new_n8156_1_;
   wire new_n8155_;
   wire new_n8154_;
   wire new_n8153_;
   wire new_n8151_;
   wire new_n8150_;
   wire new_n8149_;
   wire new_n8147_1_;
   wire new_n8146_;
   wire new_n8145_;
   wire new_n8144_1_;
   wire new_n8143_;
   wire new_n8142_;
   wire new_n8141_;
   wire new_n8140_1_;
   wire new_n8139_;
   wire new_n8135_1_;
   wire new_n8134_;
   wire new_n8133_;
   wire new_n8132_;
   wire new_n8131_;
   wire new_n8124_;
   wire new_n8123_;
   wire new_n8122_;
   wire new_n8121_1_;
   wire new_n8120_;
   wire new_n8119_;
   wire new_n8118_;
   wire new_n8117_;
   wire new_n8114_;
   wire new_n8113_;
   wire new_n8112_1_;
   wire new_n8107_1_;
   wire new_n8106_;
   wire new_n8105_;
   wire new_n8104_;
   wire new_n8103_;
   wire new_n8102_1_;
   wire new_n8100_;
   wire new_n8099_;
   wire new_n8091_;
   wire new_n8090_;
   wire new_n8084_;
   wire new_n8083_;
   wire new_n8082_;
   wire new_n8081_;
   wire new_n8080_1_;
   wire new_n8079_;
   wire new_n8078_;
   wire new_n8077_;
   wire new_n8076_;
   wire new_n8075_1_;
   wire new_n8074_;
   wire new_n8073_;
   wire new_n8072_1_;
   wire new_n8071_;
   wire new_n8068_;
   wire new_n8067_1_;
   wire new_n8066_;
   wire new_n8065_;
   wire new_n8064_1_;
   wire new_n8061_;
   wire new_n8060_;
   wire new_n8059_1_;
   wire new_n8058_;
   wire new_n8057_;
   wire new_n8056_1_;
   wire new_n8055_;
   wire new_n8054_;
   wire new_n8053_;
   wire new_n8052_;
   wire new_n8051_1_;
   wire new_n8050_;
   wire new_n8049_;
   wire new_n8048_;
   wire new_n8044_;
   wire new_n8043_;
   wire new_n8042_1_;
   wire new_n8041_;
   wire new_n8040_;
   wire new_n8035_;
   wire new_n8034_;
   wire new_n8033_1_;
   wire new_n8032_;
   wire new_n8031_;
   wire new_n8030_;
   wire new_n8029_;
   wire new_n8028_1_;
   wire new_n8027_;
   wire new_n8026_;
   wire new_n8025_;
   wire new_n8024_1_;
   wire new_n8023_;
   wire new_n8022_;
   wire new_n8021_;
   wire new_n8020_;
   wire new_n8011_;
   wire new_n8010_1_;
   wire new_n8009_;
   wire new_n8005_1_;
   wire new_n8004_;
   wire new_n8001_;
   wire new_n8000_;
   wire new_n7999_;
   wire new_n7993_;
   wire new_n7992_;
   wire new_n7991_;
   wire new_n7990_;
   wire new_n7989_1_;
   wire new_n7987_;
   wire new_n7986_;
   wire new_n7985_1_;
   wire new_n7983_;
   wire new_n7978_;
   wire new_n7977_;
   wire new_n7976_;
   wire new_n7975_1_;
   wire new_n7972_;
   wire new_n7971_;
   wire new_n7970_1_;
   wire new_n7965_;
   wire new_n7964_;
   wire new_n7963_;
   wire new_n7962_1_;
   wire new_n7961_;
   wire new_n7960_;
   wire new_n7957_;
   wire new_n7956_;
   wire new_n7955_1_;
   wire new_n7954_;
   wire new_n7953_;
   wire new_n7952_;
   wire new_n7951_;
   wire new_n7950_1_;
   wire new_n7949_;
   wire new_n7946_;
   wire new_n7945_1_;
   wire new_n7944_;
   wire new_n7943_;
   wire new_n7942_1_;
   wire new_n7941_;
   wire new_n7940_;
   wire new_n7939_;
   wire new_n7938_;
   wire new_n7937_1_;
   wire new_n7936_;
   wire new_n7935_;
   wire new_n7934_;
   wire new_n7931_;
   wire new_n7930_;
   wire new_n7929_1_;
   wire new_n7925_;
   wire new_n7924_1_;
   wire new_n7923_;
   wire new_n7922_;
   wire new_n7921_;
   wire new_n7920_1_;
   wire new_n7919_;
   wire new_n7918_;
   wire new_n7917_;
   wire new_n7916_1_;
   wire new_n7915_;
   wire new_n7914_;
   wire new_n7913_;
   wire new_n7912_;
   wire new_n7911_1_;
   wire new_n7910_;
   wire new_n7909_;
   wire new_n7908_;
   wire new_n7907_;
   wire new_n7906_1_;
   wire new_n7905_;
   wire new_n7904_;
   wire new_n7903_;
   wire new_n7902_1_;
   wire new_n7896_;
   wire new_n7895_;
   wire new_n7892_;
   wire new_n7891_;
   wire new_n7878_1_;
   wire new_n7876_;
   wire new_n7875_1_;
   wire new_n7874_;
   wire new_n7873_;
   wire new_n7872_;
   wire new_n7869_;
   wire new_n7868_;
   wire new_n7865_;
   wire new_n7864_;
   wire new_n7863_1_;
   wire new_n7862_;
   wire new_n7861_;
   wire new_n7860_;
   wire new_n7859_;
   wire new_n7858_1_;
   wire new_n7857_;
   wire new_n7856_;
   wire new_n7855_;
   wire new_n7854_;
   wire new_n7853_1_;
   wire new_n7851_;
   wire new_n7850_;
   wire new_n7849_;
   wire new_n7848_1_;
   wire new_n7847_;
   wire new_n7845_1_;
   wire new_n7844_;
   wire new_n7843_;
   wire new_n7842_;
   wire new_n7841_;
   wire new_n7840_1_;
   wire new_n7839_;
   wire new_n7838_;
   wire new_n7837_;
   wire new_n7836_;
   wire new_n7835_1_;
   wire new_n7834_;
   wire new_n7833_;
   wire new_n7832_;
   wire new_n7831_1_;
   wire new_n7830_;
   wire new_n7829_;
   wire new_n7828_;
   wire new_n7827_;
   wire new_n7826_1_;
   wire new_n7825_;
   wire new_n7824_;
   wire new_n7823_;
   wire new_n7822_1_;
   wire new_n7821_;
   wire new_n7820_;
   wire new_n7819_;
   wire new_n7818_1_;
   wire new_n7817_;
   wire new_n7816_;
   wire new_n7815_1_;
   wire new_n7814_;
   wire new_n7813_;
   wire new_n7812_;
   wire new_n7811_;
   wire new_n7810_1_;
   wire new_n7806_1_;
   wire new_n7805_;
   wire new_n7804_;
   wire new_n7798_1_;
   wire new_n7797_;
   wire new_n7796_;
   wire new_n7795_;
   wire new_n7794_;
   wire new_n7792_;
   wire new_n7791_;
   wire new_n7779_1_;
   wire new_n7775_;
   wire new_n7774_;
   wire new_n7773_1_;
   wire new_n7772_;
   wire new_n7771_;
   wire new_n7767_;
   wire new_n7766_;
   wire new_n7762_;
   wire new_n7761_;
   wire new_n7760_1_;
   wire new_n7756_1_;
   wire new_n7755_;
   wire new_n7754_;
   wire new_n7753_;
   wire new_n7752_;
   wire new_n7747_;
   wire new_n7744_;
   wire new_n7741_1_;
   wire new_n7740_;
   wire new_n7739_;
   wire new_n7738_;
   wire new_n7736_;
   wire new_n7735_;
   wire new_n7734_;
   wire new_n7733_;
   wire new_n7732_1_;
   wire new_n7731_;
   wire new_n7730_;
   wire new_n7721_;
   wire new_n7720_;
   wire new_n7719_1_;
   wire new_n7718_;
   wire new_n7717_;
   wire new_n7716_;
   wire new_n7715_;
   wire new_n7714_1_;
   wire new_n7713_;
   wire new_n7712_;
   wire new_n7711_;
   wire new_n7710_;
   wire new_n7709_1_;
   wire new_n7708_;
   wire new_n7702_;
   wire new_n7701_;
   wire new_n7700_1_;
   wire new_n7699_;
   wire new_n7698_;
   wire new_n7697_;
   wire new_n7696_;
   wire new_n7695_1_;
   wire new_n7694_;
   wire new_n7693_;
   wire new_n7692_;
   wire new_n7691_1_;
   wire new_n7690_;
   wire new_n7689_;
   wire new_n7688_;
   wire new_n7687_;
   wire new_n7686_1_;
   wire new_n7685_;
   wire new_n7684_;
   wire new_n7683_;
   wire new_n7682_;
   wire new_n7681_1_;
   wire new_n7680_;
   wire new_n7679_;
   wire new_n7678_;
   wire new_n7677_;
   wire new_n7676_1_;
   wire new_n7675_;
   wire new_n7674_;
   wire new_n7669_;
   wire new_n7668_;
   wire new_n7667_;
   wire new_n7666_1_;
   wire new_n7665_;
   wire new_n7662_;
   wire new_n7661_1_;
   wire new_n7657_;
   wire new_n7656_;
   wire new_n7655_;
   wire new_n7652_;
   wire new_n7651_;
   wire new_n7650_;
   wire new_n7649_1_;
   wire new_n7648_;
   wire new_n7647_;
   wire new_n7646_;
   wire new_n7645_;
   wire new_n7644_1_;
   wire new_n7643_;
   wire new_n7633_;
   wire new_n7632_;
   wire new_n7631_1_;
   wire new_n7630_;
   wire new_n7629_;
   wire new_n7626_1_;
   wire new_n7625_;
   wire new_n7624_;
   wire new_n7623_;
   wire new_n7622_1_;
   wire new_n7621_;
   wire new_n7620_;
   wire new_n7619_;
   wire new_n7618_1_;
   wire new_n7617_;
   wire new_n7616_;
   wire new_n7615_;
   wire new_n7614_;
   wire new_n7613_1_;
   wire new_n7612_;
   wire new_n7609_;
   wire new_n7608_1_;
   wire new_n7605_;
   wire new_n7604_1_;
   wire new_n7602_;
   wire new_n7597_;
   wire new_n7596_1_;
   wire new_n7595_;
   wire new_n7594_;
   wire new_n7593_;
   wire new_n7590_;
   wire new_n7589_;
   wire new_n7588_;
   wire new_n7587_;
   wire new_n7586_1_;
   wire new_n7585_;
   wire new_n7584_;
   wire new_n7583_;
   wire new_n7582_;
   wire new_n7581_1_;
   wire new_n7580_;
   wire new_n7579_;
   wire new_n7578_;
   wire new_n7577_1_;
   wire new_n7576_;
   wire new_n7575_;
   wire new_n7574_;
   wire new_n7573_;
   wire new_n7572_1_;
   wire new_n7571_;
   wire new_n7570_;
   wire new_n7569_;
   wire new_n7568_;
   wire new_n7567_1_;
   wire new_n7566_;
   wire new_n7565_;
   wire new_n7564_;
   wire new_n7563_1_;
   wire new_n7562_;
   wire new_n7561_;
   wire new_n7560_;
   wire new_n7559_;
   wire new_n7558_1_;
   wire new_n7557_;
   wire new_n7556_;
   wire new_n7555_;
   wire new_n7554_;
   wire new_n7553_1_;
   wire new_n7552_;
   wire new_n7547_;
   wire new_n7545_;
   wire new_n7544_;
   wire new_n7543_1_;
   wire new_n7542_;
   wire new_n7541_;
   wire new_n7540_;
   wire new_n7538_;
   wire new_n7537_;
   wire new_n7533_;
   wire new_n7532_;
   wire new_n7531_;
   wire new_n7530_1_;
   wire new_n7529_;
   wire new_n7527_1_;
   wire new_n7526_;
   wire new_n7525_;
   wire new_n7523_;
   wire new_n7522_1_;
   wire new_n7521_;
   wire new_n7516_;
   wire new_n7515_;
   wire new_n7513_1_;
   wire new_n7512_;
   wire new_n7511_;
   wire new_n7510_;
   wire new_n7509_1_;
   wire new_n7508_;
   wire new_n7504_;
   wire new_n7503_;
   wire new_n7502_;
   wire new_n7501_1_;
   wire new_n7500_;
   wire new_n7499_;
   wire new_n7497_;
   wire new_n7496_1_;
   wire new_n7495_;
   wire new_n7494_;
   wire new_n7493_;
   wire new_n7492_1_;
   wire new_n7486_;
   wire new_n7485_;
   wire new_n7484_;
   wire new_n7483_;
   wire new_n7482_1_;
   wire new_n7472_;
   wire new_n7471_;
   wire new_n7467_;
   wire new_n7466_;
   wire new_n7465_;
   wire new_n7461_;
   wire new_n7460_;
   wire new_n7459_1_;
   wire new_n7452_;
   wire new_n7451_;
   wire new_n7450_1_;
   wire new_n7449_;
   wire new_n7448_;
   wire new_n7447_;
   wire new_n7446_1_;
   wire new_n7445_;
   wire new_n7444_;
   wire new_n7443_;
   wire new_n7442_1_;
   wire new_n7437_1_;
   wire new_n7436_;
   wire new_n7435_;
   wire new_n7430_;
   wire new_n7429_;
   wire new_n7428_;
   wire new_n7427_1_;
   wire new_n7424_;
   wire new_n7423_;
   wire new_n7422_1_;
   wire new_n7418_;
   wire new_n7417_1_;
   wire new_n7416_;
   wire new_n7415_;
   wire new_n7414_;
   wire new_n7413_1_;
   wire new_n7412_;
   wire new_n7411_;
   wire new_n7408_1_;
   wire new_n7407_;
   wire new_n7404_1_;
   wire new_n7403_;
   wire new_n7401_;
   wire new_n7400_1_;
   wire new_n7399_;
   wire new_n7398_;
   wire new_n7397_;
   wire new_n7396_;
   wire new_n7395_1_;
   wire new_n7394_;
   wire new_n7393_;
   wire new_n7392_;
   wire new_n7391_1_;
   wire new_n7390_;
   wire new_n7389_;
   wire new_n7388_;
   wire new_n7387_;
   wire new_n7386_1_;
   wire new_n7385_;
   wire new_n7384_;
   wire new_n7383_;
   wire new_n7382_;
   wire new_n7381_1_;
   wire new_n7380_;
   wire new_n7379_;
   wire new_n7378_;
   wire new_n7377_;
   wire new_n7376_1_;
   wire new_n7375_;
   wire new_n7374_;
   wire new_n7373_;
   wire new_n7372_1_;
   wire new_n7371_;
   wire new_n7370_;
   wire new_n7369_;
   wire new_n7368_1_;
   wire new_n7367_;
   wire new_n7366_;
   wire new_n7365_;
   wire new_n7364_;
   wire new_n7363_1_;
   wire new_n7362_;
   wire new_n7361_;
   wire new_n7360_;
   wire new_n7359_1_;
   wire new_n7358_;
   wire new_n7357_;
   wire new_n7356_;
   wire new_n7355_;
   wire new_n7354_1_;
   wire new_n7352_;
   wire new_n7351_;
   wire new_n7350_;
   wire new_n7346_;
   wire new_n7345_;
   wire new_n7344_1_;
   wire new_n7343_;
   wire new_n7342_;
   wire new_n7341_;
   wire new_n7340_1_;
   wire new_n7339_;
   wire new_n7337_;
   wire new_n7336_;
   wire new_n7335_1_;
   wire new_n7334_;
   wire new_n7333_;
   wire new_n7329_;
   wire new_n7328_;
   wire new_n7326_1_;
   wire new_n7325_;
   wire new_n7323_;
   wire new_n7322_;
   wire new_n7321_1_;
   wire new_n7320_;
   wire new_n7319_;
   wire new_n7312_1_;
   wire new_n7311_;
   wire new_n7310_;
   wire new_n7309_;
   wire new_n7306_;
   wire new_n7305_;
   wire new_n7304_;
   wire new_n7303_;
   wire new_n7302_1_;
   wire new_n7301_;
   wire new_n7300_;
   wire new_n7299_;
   wire new_n7298_;
   wire new_n7297_1_;
   wire new_n7296_;
   wire new_n7295_;
   wire new_n7294_;
   wire new_n7292_1_;
   wire new_n7291_;
   wire new_n7290_;
   wire new_n7289_;
   wire new_n7288_1_;
   wire new_n7287_;
   wire new_n7285_;
   wire new_n7284_1_;
   wire new_n7283_;
   wire new_n7282_;
   wire new_n7279_;
   wire new_n7278_;
   wire new_n7277_;
   wire new_n7276_;
   wire new_n7275_1_;
   wire new_n7274_;
   wire new_n7273_;
   wire new_n7272_;
   wire new_n7271_;
   wire new_n7270_1_;
   wire new_n7269_;
   wire new_n7268_;
   wire new_n7265_1_;
   wire new_n7264_;
   wire new_n7262_;
   wire new_n7258_;
   wire new_n7257_;
   wire new_n7256_1_;
   wire new_n7255_;
   wire new_n7254_;
   wire new_n7253_;
   wire new_n7252_1_;
   wire new_n7251_;
   wire new_n7250_;
   wire new_n7249_1_;
   wire new_n7248_;
   wire new_n7239_;
   wire new_n7236_;
   wire new_n7235_1_;
   wire new_n7234_;
   wire new_n7233_;
   wire new_n7232_;
   wire new_n7230_1_;
   wire new_n7229_;
   wire new_n7228_;
   wire new_n7227_;
   wire new_n7225_;
   wire new_n7224_;
   wire new_n7223_;
   wire new_n7222_;
   wire new_n7221_1_;
   wire new_n7220_;
   wire new_n7219_;
   wire new_n7218_;
   wire new_n7216_1_;
   wire new_n7215_;
   wire new_n7214_;
   wire new_n7213_;
   wire new_n7211_;
   wire new_n7210_;
   wire new_n7209_;
   wire new_n7208_;
   wire new_n7207_1_;
   wire new_n7206_;
   wire new_n7205_;
   wire new_n7204_;
   wire new_n7203_1_;
   wire new_n7202_;
   wire new_n7201_;
   wire new_n7200_;
   wire new_n7199_1_;
   wire new_n7198_;
   wire new_n7197_;
   wire new_n7196_;
   wire new_n7195_;
   wire new_n7194_1_;
   wire new_n7193_;
   wire new_n7192_;
   wire new_n7191_;
   wire new_n7190_1_;
   wire new_n7189_;
   wire new_n7188_;
   wire new_n7187_;
   wire new_n7186_;
   wire new_n7184_;
   wire new_n7183_;
   wire new_n7182_1_;
   wire new_n7181_;
   wire new_n7179_;
   wire new_n7178_;
   wire new_n7177_1_;
   wire new_n7175_;
   wire new_n7174_;
   wire new_n7173_;
   wire new_n7172_1_;
   wire new_n7171_;
   wire new_n7170_;
   wire new_n7169_;
   wire new_n7168_;
   wire new_n7167_1_;
   wire new_n7166_;
   wire new_n7165_;
   wire new_n7164_1_;
   wire new_n7163_;
   wire new_n7162_;
   wire new_n7161_;
   wire new_n7160_1_;
   wire new_n7159_;
   wire new_n7158_;
   wire new_n7157_;
   wire new_n7156_;
   wire new_n7155_1_;
   wire new_n7154_;
   wire new_n7153_;
   wire new_n7152_;
   wire new_n7151_1_;
   wire new_n7148_;
   wire new_n7137_;
   wire new_n7136_;
   wire new_n7135_;
   wire new_n7134_;
   wire new_n7133_1_;
   wire new_n7132_;
   wire new_n7131_;
   wire new_n7130_;
   wire new_n7129_;
   wire new_n7128_1_;
   wire new_n7127_;
   wire new_n7126_;
   wire new_n7125_1_;
   wire new_n7124_;
   wire new_n7123_;
   wire new_n7122_;
   wire new_n7121_;
   wire new_n7120_1_;
   wire new_n7119_;
   wire new_n7118_;
   wire new_n7117_;
   wire new_n7116_1_;
   wire new_n7115_;
   wire new_n7114_;
   wire new_n7113_;
   wire new_n7111_1_;
   wire new_n7110_;
   wire new_n7109_;
   wire new_n7108_;
   wire new_n7107_1_;
   wire new_n7106_;
   wire new_n7105_;
   wire new_n7104_;
   wire new_n7103_;
   wire new_n7102_1_;
   wire new_n7101_;
   wire new_n7100_;
   wire new_n7099_;
   wire new_n7098_1_;
   wire new_n7097_;
   wire new_n7093_1_;
   wire new_n7092_;
   wire new_n7091_;
   wire new_n7090_;
   wire new_n7089_1_;
   wire new_n7088_;
   wire new_n7087_;
   wire new_n7086_;
   wire new_n7085_1_;
   wire new_n7084_;
   wire new_n7083_;
   wire new_n7082_1_;
   wire new_n7081_;
   wire new_n7080_;
   wire new_n7079_;
   wire new_n7078_;
   wire new_n7077_1_;
   wire new_n7076_;
   wire new_n7075_;
   wire new_n7074_;
   wire new_n7073_;
   wire new_n7072_1_;
   wire new_n7071_;
   wire new_n7070_;
   wire new_n7069_;
   wire new_n7068_;
   wire new_n7067_1_;
   wire new_n7066_;
   wire new_n7065_;
   wire new_n7064_;
   wire new_n7063_;
   wire new_n7062_1_;
   wire new_n7061_;
   wire new_n7060_;
   wire new_n7059_;
   wire new_n7058_1_;
   wire new_n7057_;
   wire new_n7056_;
   wire new_n7055_;
   wire new_n7054_;
   wire new_n7053_1_;
   wire new_n7052_;
   wire new_n7051_;
   wire new_n7050_;
   wire new_n7049_1_;
   wire new_n7048_;
   wire new_n7047_;
   wire new_n7046_;
   wire new_n7045_1_;
   wire new_n7044_;
   wire new_n7043_;
   wire new_n7042_;
   wire new_n7035_;
   wire new_n7034_;
   wire new_n7029_;
   wire new_n7028_;
   wire new_n7027_1_;
   wire new_n7026_;
   wire new_n7025_;
   wire new_n7024_;
   wire new_n7023_1_;
   wire new_n7022_;
   wire new_n7021_;
   wire new_n7020_;
   wire new_n7019_;
   wire new_n7018_1_;
   wire new_n7017_;
   wire new_n7014_;
   wire new_n7013_1_;
   wire new_n7012_;
   wire new_n7011_;
   wire new_n7010_;
   wire new_n7009_1_;
   wire new_n7008_;
   wire new_n7007_;
   wire new_n7006_;
   wire new_n7005_1_;
   wire new_n7004_;
   wire new_n7003_;
   wire new_n7002_;
   wire new_n7001_;
   wire new_n7000_1_;
   wire new_n6999_;
   wire new_n6998_;
   wire new_n6997_;
   wire new_n6996_;
   wire new_n6995_1_;
   wire new_n6994_;
   wire new_n6993_;
   wire new_n6992_;
   wire new_n6991_;
   wire new_n6990_1_;
   wire new_n6989_;
   wire new_n6988_;
   wire new_n6987_;
   wire new_n6986_1_;
   wire new_n6985_;
   wire new_n6984_;
   wire new_n6983_;
   wire new_n6982_1_;
   wire new_n6981_;
   wire new_n6980_;
   wire new_n6979_;
   wire new_n6978_;
   wire new_n6977_1_;
   wire new_n6976_;
   wire new_n6975_;
   wire new_n6974_1_;
   wire new_n6973_;
   wire new_n6972_;
   wire new_n6971_;
   wire new_n6970_;
   wire new_n6969_1_;
   wire new_n6968_;
   wire new_n6967_;
   wire new_n6966_;
   wire new_n6965_;
   wire new_n6963_;
   wire new_n6961_;
   wire new_n6960_1_;
   wire new_n6959_;
   wire new_n6957_1_;
   wire new_n6956_;
   wire new_n6955_;
   wire new_n6954_;
   wire new_n6953_;
   wire new_n6952_1_;
   wire new_n6951_;
   wire new_n6950_;
   wire new_n6949_;
   wire new_n6948_;
   wire new_n6947_1_;
   wire new_n6946_;
   wire new_n6945_;
   wire new_n6944_;
   wire new_n6943_1_;
   wire new_n6942_;
   wire new_n6941_;
   wire new_n6940_;
   wire new_n6939_;
   wire new_n6937_;
   wire new_n6936_;
   wire new_n6935_;
   wire new_n6934_1_;
   wire new_n6933_;
   wire new_n6932_;
   wire new_n6920_;
   wire new_n6919_1_;
   wire new_n6918_;
   wire new_n6917_;
   wire new_n6916_;
   wire new_n6915_1_;
   wire new_n6914_;
   wire new_n6913_;
   wire new_n6912_;
   wire new_n6911_;
   wire new_n6910_1_;
   wire new_n6909_;
   wire new_n6907_;
   wire new_n6906_1_;
   wire new_n6905_;
   wire new_n6904_;
   wire new_n6903_;
   wire new_n6902_1_;
   wire new_n6901_;
   wire new_n6900_;
   wire new_n6899_1_;
   wire new_n6898_;
   wire new_n6897_;
   wire new_n6896_;
   wire new_n6895_1_;
   wire new_n6894_;
   wire new_n6893_;
   wire new_n6892_;
   wire new_n6891_;
   wire new_n6890_1_;
   wire new_n6889_;
   wire new_n6888_;
   wire new_n6887_;
   wire new_n6886_1_;
   wire new_n6882_;
   wire new_n6881_1_;
   wire new_n6880_;
   wire new_n6879_;
   wire new_n6878_;
   wire new_n6877_;
   wire new_n6876_1_;
   wire new_n6875_;
   wire new_n6874_;
   wire new_n6873_;
   wire new_n6872_1_;
   wire new_n6871_;
   wire new_n6870_;
   wire new_n6869_;
   wire new_n6868_;
   wire new_n6867_1_;
   wire new_n6866_;
   wire new_n6865_;
   wire new_n6864_;
   wire new_n6863_1_;
   wire new_n6862_;
   wire new_n6861_;
   wire new_n6860_1_;
   wire new_n6859_;
   wire new_n6858_;
   wire new_n6857_;
   wire new_n6856_;
   wire new_n6855_1_;
   wire new_n6854_;
   wire new_n6853_;
   wire new_n6852_;
   wire new_n6851_;
   wire new_n6850_1_;
   wire new_n6849_;
   wire new_n6848_;
   wire new_n6847_;
   wire new_n6846_;
   wire new_n6845_1_;
   wire new_n6844_;
   wire new_n6843_;
   wire new_n6842_;
   wire new_n6841_;
   wire new_n6840_1_;
   wire new_n6839_;
   wire new_n6838_;
   wire new_n6837_;
   wire new_n6836_1_;
   wire new_n6835_;
   wire new_n6834_;
   wire new_n6833_;
   wire new_n6832_;
   wire new_n6831_1_;
   wire new_n6830_;
   wire new_n6829_;
   wire new_n6828_;
   wire new_n6827_;
   wire new_n6826_1_;
   wire new_n6825_;
   wire new_n6823_;
   wire new_n6822_1_;
   wire new_n6821_;
   wire new_n6820_;
   wire new_n6819_;
   wire new_n6815_;
   wire new_n6814_;
   wire new_n6813_1_;
   wire new_n6812_;
   wire new_n6811_;
   wire new_n6810_;
   wire new_n6809_1_;
   wire new_n6808_;
   wire new_n6807_;
   wire new_n6806_1_;
   wire new_n6805_;
   wire new_n6804_;
   wire new_n6803_;
   wire new_n6802_;
   wire new_n6801_1_;
   wire new_n6800_;
   wire new_n6799_;
   wire new_n6798_;
   wire new_n6797_;
   wire new_n6796_1_;
   wire new_n6795_;
   wire new_n6794_;
   wire new_n6793_1_;
   wire new_n6792_;
   wire new_n6791_;
   wire new_n6790_;
   wire new_n6789_;
   wire new_n6788_1_;
   wire new_n6787_;
   wire new_n6786_;
   wire new_n6785_;
   wire new_n6784_;
   wire new_n6783_1_;
   wire new_n6782_;
   wire new_n6781_;
   wire new_n6780_;
   wire new_n6779_1_;
   wire new_n6778_;
   wire new_n6777_;
   wire new_n6776_;
   wire new_n6775_;
   wire new_n6774_1_;
   wire new_n6773_;
   wire new_n6772_;
   wire new_n6771_;
   wire new_n6770_1_;
   wire new_n6769_;
   wire new_n6768_;
   wire new_n6767_;
   wire new_n6766_;
   wire new_n6765_1_;
   wire new_n6764_;
   wire new_n6763_;
   wire new_n6762_;
   wire new_n6761_1_;
   wire new_n6760_;
   wire new_n6759_;
   wire new_n6756_1_;
   wire new_n6755_;
   wire new_n6754_;
   wire new_n6752_1_;
   wire new_n6751_;
   wire new_n6750_;
   wire new_n6749_1_;
   wire new_n6748_;
   wire new_n6747_;
   wire new_n6746_1_;
   wire new_n6745_;
   wire new_n6744_;
   wire new_n6743_;
   wire new_n6742_;
   wire new_n6741_1_;
   wire new_n12336_;
   wire new_n12332_;
   wire new_n12331_;
   wire new_n12330_;
   wire new_n12329_;
   wire new_n12328_;
   wire new_n12327_;
   wire new_n12326_;
   wire new_n12325_;
   wire new_n12324_;
   wire new_n12321_;
   wire new_n12317_;
   wire new_n12316_;
   wire new_n12311_;
   wire new_n12309_;
   wire new_n12308_;
   wire new_n12306_;
   wire new_n12305_;
   wire new_n12304_;
   wire new_n12303_;
   wire new_n12302_;
   wire new_n12301_;
   wire new_n12300_;
   wire new_n12299_;
   wire new_n12298_;
   wire new_n12296_;
   wire new_n12295_;
   wire new_n12294_;
   wire new_n12293_;
   wire new_n12291_;
   wire new_n12290_;
   wire new_n12289_;
   wire new_n12287_;
   wire new_n12286_;
   wire new_n12283_;
   wire new_n12282_;
   wire new_n12281_;
   wire new_n12280_;
   wire new_n12279_;
   wire new_n12278_;
   wire new_n12277_;
   wire new_n12276_;
   wire new_n12275_;
   wire new_n12274_;
   wire new_n12273_;
   wire new_n12272_;
   wire new_n12271_;
   wire new_n12269_;
   wire new_n12266_;
   wire new_n12249_;
   wire new_n12246_;
   wire new_n12245_;
   wire new_n12244_;
   wire new_n12243_;
   wire new_n12242_;
   wire new_n12241_;
   wire new_n12240_;
   wire new_n12239_;
   wire new_n12238_;
   wire new_n12236_;
   wire new_n12235_;
   wire new_n12230_;
   wire new_n12227_;
   wire new_n12218_;
   wire new_n12217_;
   wire new_n12216_;
   wire new_n12215_;
   wire new_n12214_;
   wire new_n12213_;
   wire new_n12212_;
   wire new_n12211_;
   wire new_n12210_;
   wire new_n12209_;
   wire new_n12205_;
   wire new_n12204_;
   wire new_n12202_;
   wire new_n12201_;
   wire new_n12200_;
   wire new_n12199_;
   wire new_n12196_;
   wire new_n12195_;
   wire new_n12190_;
   wire new_n12188_;
   wire new_n12185_;
   wire new_n12184_;
   wire new_n12177_;
   wire new_n12176_;
   wire new_n12175_;
   wire new_n12174_;
   wire new_n12172_;
   wire new_n12170_;
   wire new_n12166_;
   wire new_n12165_;
   wire new_n12164_;
   wire new_n12163_;
   wire new_n12162_;
   wire new_n12155_;
   wire new_n12148_;
   wire new_n12145_;
   wire new_n12141_;
   wire new_n12140_;
   wire new_n12139_;
   wire new_n12138_;
   wire new_n12137_;
   wire new_n12136_;
   wire new_n12135_;
   wire new_n12134_;
   wire new_n12133_;
   wire new_n12131_;
   wire new_n12130_;
   wire new_n12129_;
   wire new_n12128_;
   wire new_n12127_;
   wire new_n12126_;
   wire new_n12125_;
   wire new_n12124_;
   wire new_n12123_;
   wire new_n12122_;
   wire new_n12121_;
   wire new_n12120_;
   wire new_n12119_;
   wire new_n12118_;
   wire new_n12114_;
   wire new_n12113_;
   wire new_n12112_;
   wire new_n12111_;
   wire new_n12110_;
   wire new_n12109_;
   wire new_n12103_;
   wire new_n12097_;
   wire new_n12096_;
   wire new_n12091_;
   wire new_n12090_;
   wire new_n12088_;
   wire new_n12087_;
   wire new_n12079_;
   wire new_n12078_;
   wire new_n12076_;
   wire new_n12075_;
   wire new_n12074_;
   wire new_n12073_;
   wire new_n12072_;
   wire new_n12071_;
   wire new_n12070_;
   wire new_n12069_;
   wire new_n12068_;
   wire new_n12065_;
   wire new_n12061_;
   wire new_n12057_;
   wire new_n12056_;
   wire new_n12053_;
   wire new_n12052_;
   wire new_n12051_;
   wire new_n12050_;
   wire new_n12049_;
   wire new_n12048_;
   wire new_n12047_;
   wire new_n12046_;
   wire new_n12045_;
   wire new_n12044_;
   wire new_n12043_;
   wire new_n12042_;
   wire new_n12041_;
   wire new_n12040_;
   wire new_n12039_;
   wire new_n12038_;
   wire new_n12037_;
   wire new_n12036_;
   wire new_n12035_;
   wire new_n12031_;
   wire new_n12030_;
   wire new_n12020_;
   wire new_n12018_;
   wire new_n12017_;
   wire new_n12008_;
   wire new_n12007_;
   wire new_n12006_;
   wire new_n12005_;
   wire new_n12004_;
   wire new_n12000_;
   wire new_n11999_;
   wire new_n11998_;
   wire new_n11997_;
   wire new_n11996_;
   wire new_n11995_;
   wire new_n11994_;
   wire new_n11993_;
   wire new_n11992_;
   wire new_n11991_;
   wire new_n11990_;
   wire new_n11989_;
   wire new_n11987_;
   wire new_n11982_;
   wire new_n11981_;
   wire new_n11979_;
   wire new_n11978_;
   wire new_n11962_;
   wire new_n11957_;
   wire new_n11953_;
   wire new_n11952_;
   wire new_n11948_;
   wire new_n11941_;
   wire new_n11940_;
   wire new_n11939_;
   wire new_n11938_;
   wire new_n11937_;
   wire new_n11936_;
   wire new_n11935_;
   wire new_n11934_;
   wire new_n11933_;
   wire new_n11931_;
   wire new_n11930_;
   wire new_n11928_;
   wire new_n11927_;
   wire new_n11924_;
   wire new_n11922_;
   wire new_n11912_;
   wire new_n11911_;
   wire new_n11910_;
   wire new_n11909_;
   wire new_n11908_;
   wire new_n11907_;
   wire new_n11906_;
   wire new_n11905_;
   wire new_n11904_;
   wire new_n11901_;
   wire new_n11898_;
   wire new_n11895_;
   wire new_n11893_;
   wire new_n11892_;
   wire new_n11884_;
   wire new_n11883_;
   wire new_n11881_;
   wire new_n11868_;
   wire new_n11867_;
   wire new_n11856_;
   wire new_n11855_;
   wire new_n11852_;
   wire new_n11851_;
   wire new_n11847_;
   wire new_n11846_;
   wire new_n11845_;
   wire new_n11844_;
   wire new_n11843_;
   wire new_n11842_;
   wire new_n11841_;
   wire new_n11840_;
   wire new_n11839_;
   wire new_n11832_;
   wire new_n11831_;
   wire new_n11829_;
   wire new_n11823_;
   wire new_n11820_;
   wire new_n11816_;
   wire new_n11815_;
   wire new_n11813_;
   wire new_n11812_;
   wire new_n11805_;
   wire new_n11803_;
   wire new_n11802_;
   wire new_n11787_;
   wire new_n11785_;
   wire new_n11784_;
   wire new_n11780_;
   wire new_n11776_;
   wire new_n11775_;
   wire new_n11772_;
   wire new_n11764_;
   wire new_n11763_;
   wire new_n11761_;
   wire new_n11760_;
   wire new_n11759_;
   wire new_n11758_;
   wire new_n11757_;
   wire new_n11755_;
   wire new_n11749_;
   wire new_n11744_;
   wire new_n11743_;
   wire new_n11742_;
   wire new_n11741_;
   wire new_n11739_;
   wire new_n11738_;
   wire new_n11736_;
   wire new_n11732_;
   wire new_n11731_;
   wire new_n11730_;
   wire new_n11729_;
   wire new_n11728_;
   wire new_n11727_;
   wire new_n11726_;
   wire new_n11725_;
   wire new_n11724_;
   wire new_n11723_;
   wire new_n11722_;
   wire new_n11721_;
   wire new_n11720_;
   wire new_n11716_;
   wire new_n11715_;
   wire new_n11709_;
   wire new_n11708_;
   wire new_n11705_;
   wire new_n11700_;
   wire new_n11699_;
   wire new_n11698_;
   wire new_n11697_;
   wire new_n11696_;
   wire new_n11695_;
   wire new_n11694_;
   wire new_n11693_;
   wire new_n11692_;
   wire new_n11686_;
   wire new_n11683_;
   wire new_n11680_;
   wire new_n11679_;
   wire new_n11678_;
   wire new_n11676_;
   wire new_n11675_;
   wire new_n11671_;
   wire new_n11663_;
   wire new_n11662_;
   wire new_n11657_;
   wire new_n11656_;
   wire new_n11653_;
   wire new_n11651_;
   wire new_n11646_;
   wire new_n11640_;
   wire new_n11639_;
   wire new_n11638_;
   wire new_n11637_;
   wire new_n11636_;
   wire new_n11635_;
   wire new_n11634_;
   wire new_n11633_;
   wire new_n11632_;
   wire new_n11631_;
   wire new_n11630_;
   wire new_n11629_;
   wire new_n11628_;
   wire new_n11627_;
   wire new_n11625_;
   wire new_n11624_;
   wire new_n11613_;
   wire new_n11612_;
   wire new_n11611_;
   wire new_n11610_;
   wire new_n11609_;
   wire new_n11608_;
   wire new_n11607_;
   wire new_n11606_;
   wire new_n11605_;
   wire new_n11604_;
   wire new_n11601_;
   wire new_n11600_;
   wire new_n11599_;
   wire new_n11598_;
   wire new_n11593_;
   wire new_n11592_;
   wire new_n11590_;
   wire new_n11589_;
   wire new_n11584_;
   wire new_n11583_;
   wire new_n11582_;
   wire new_n11581_;
   wire new_n11578_;
   wire new_n11576_;
   wire new_n11575_;
   wire new_n11574_;
   wire new_n11573_;
   wire new_n11568_;
   wire new_n11567_;
   wire new_n11564_;
   wire new_n11563_;
   wire new_n11562_;
   wire new_n11561_;
   wire new_n11560_;
   wire new_n11559_;
   wire new_n11558_;
   wire new_n11557_;
   wire new_n11556_;
   wire new_n11555_;
   wire new_n11554_;
   wire new_n11553_;
   wire new_n11552_;
   wire new_n11551_;
   wire new_n11550_;
   wire new_n11535_;
   wire new_n11534_;
   wire new_n11527_;
   wire new_n11525_;
   wire new_n11524_;
   wire new_n11513_;
   wire new_n11512_;
   wire new_n11509_;
   wire new_n11508_;
   wire new_n11507_;
   wire new_n11506_;
   wire new_n11505_;
   wire new_n11504_;
   wire new_n11503_;
   wire new_n11502_;
   wire new_n11501_;
   wire new_n11499_;
   wire new_n11498_;
   wire new_n11494_;
   wire new_n11493_;
   wire new_n11492_;
   wire new_n11489_;
   wire new_n11488_;
   wire new_n11485_;
   wire new_n11484_;
   wire new_n11481_;
   wire new_n11475_;
   wire new_n11470_;
   wire new_n11469_;
   wire new_n11468_;
   wire new_n11467_;
   wire new_n11466_;
   wire new_n11465_;
   wire new_n11464_;
   wire new_n11463_;
   wire new_n11462_;
   wire new_n11461_;
   wire new_n11459_;
   wire new_n11458_;
   wire new_n11456_;
   wire new_n11455_;
   wire new_n11449_;
   wire new_n11448_;
   wire new_n11436_;
   wire new_n11435_;
   wire new_n11434_;
   wire new_n11433_;
   wire new_n11432_;
   wire new_n11431_;
   wire new_n11430_;
   wire new_n11429_;
   wire new_n11428_;
   wire new_n11422_;
   wire new_n11421_;
   wire new_n11419_;
   wire new_n11418_;
   wire new_n11417_;
   wire new_n11416_;
   wire new_n11409_;
   wire new_n11408_;
   wire new_n11406_;
   wire new_n11405_;
   wire new_n11404_;
   wire new_n11402_;
   wire new_n11395_;
   wire new_n11394_;
   wire new_n11389_;
   wire new_n11388_;
   wire new_n11382_;
   wire new_n11381_;
   wire new_n11377_;
   wire new_n11374_;
   wire new_n11367_;
   wire new_n11364_;
   wire new_n11363_;
   wire new_n11360_;
   wire new_n11359_;
   wire new_n11358_;
   wire new_n11357_;
   wire new_n11356_;
   wire new_n11355_;
   wire new_n11354_;
   wire new_n11353_;
   wire new_n11350_;
   wire new_n11349_;
   wire new_n11345_;
   wire new_n11344_;
   wire new_n11337_;
   wire new_n11336_;
   wire new_n11334_;
   wire new_n11333_;
   wire new_n11332_;
   wire new_n11330_;
   wire new_n11329_;
   wire new_n11328_;
   wire new_n11327_;
   wire new_n11326_;
   wire new_n11325_;
   wire new_n11324_;
   wire new_n11323_;
   wire new_n11322_;
   wire new_n11317_;
   wire new_n11316_;
   wire new_n11315_;
   wire new_n11314_;
   wire new_n11313_;
   wire new_n11312_;
   wire new_n11311_;
   wire new_n11310_;
   wire new_n11309_;
   wire new_n11308_;
   wire new_n11301_;
   wire new_n11298_;
   wire new_n11297_;
   wire new_n11296_;
   wire new_n11295_;
   wire new_n11294_;
   wire new_n11293_;
   wire new_n11292_;
   wire new_n11291_;
   wire new_n11290_;
   wire new_n11289_;
   wire new_n11288_;
   wire new_n11287_;
   wire new_n11286_;
   wire new_n11285_;
   wire new_n11282_;
   wire new_n11280_;
   wire new_n11279_;
   wire new_n11271_;
   wire new_n11270_;
   wire new_n11267_;
   wire new_n11266_;
   wire new_n11265_;
   wire new_n11264_;
   wire new_n11263_;
   wire new_n11262_;
   wire new_n11261_;
   wire new_n11260_;
   wire new_n11259_;
   wire new_n11257_;
   wire new_n11256_;
   wire new_n11255_;
   wire new_n11254_;
   wire new_n11253_;
   wire new_n11252_;
   wire new_n11251_;
   wire new_n11250_;
   wire new_n11249_;
   wire new_n11248_;
   wire new_n11247_;
   wire new_n11246_;
   wire new_n11244_;
   wire new_n11243_;
   wire new_n11242_;
   wire new_n11233_;
   wire new_n11232_;
   wire new_n11227_;
   wire new_n11225_;
   wire new_n11221_;
   wire new_n11220_;
   wire new_n11214_;
   wire new_n11213_;
   wire new_n11210_;
   wire new_n11208_;
   wire new_n11207_;
   wire new_n11206_;
   wire new_n11205_;
   wire new_n11202_;
   wire new_n11201_;
   wire new_n11199_;
   wire new_n11198_;
   wire new_n11197_;
   wire new_n11195_;
   wire new_n11194_;
   wire new_n11193_;
   wire new_n11192_;
   wire new_n11191_;
   wire new_n11190_;
   wire new_n11189_;
   wire new_n11188_;
   wire new_n11187_;
   wire new_n11186_;
   wire new_n11185_;
   wire new_n11184_;
   wire new_n11183_;
   wire new_n11182_;
   wire new_n11176_;
   wire new_n11175_;
   wire new_n11169_;
   wire new_n11168_;
   wire new_n11167_;
   wire new_n11166_;
   wire new_n11163_;
   wire new_n11160_;
   wire new_n11155_;
   wire new_n11154_;
   wire new_n11148_;
   wire new_n11147_;
   wire new_n11146_;
   wire new_n11145_;
   wire new_n11141_;
   wire new_n11140_;
   wire new_n11134_;
   wire new_n11130_;
   wire new_n11129_;
   wire new_n11123_;
   wire new_n11122_;
   wire new_n11121_;
   wire new_n11118_;
   wire new_n11117_;
   wire new_n11113_;
   wire new_n11112_;
   wire new_n11111_;
   wire new_n11110_;
   wire new_n11109_;
   wire new_n11108_;
   wire new_n11107_;
   wire new_n11106_;
   wire new_n11105_;
   wire new_n11100_;
   wire new_n11090_;
   wire new_n11087_;
   wire new_n11086_;
   wire new_n11085_;
   wire new_n11084_;
   wire new_n11077_;
   wire new_n11076_;
   wire new_n11074_;
   wire new_n11073_;
   wire new_n11067_;
   wire new_n11064_;
   wire new_n11063_;
   wire new_n11062_;
   wire new_n11061_;
   wire new_n11060_;
   wire new_n11059_;
   wire new_n11058_;
   wire new_n11057_;
   wire new_n11056_;
   wire new_n11052_;
   wire new_n11047_;
   wire new_n11046_;
   wire new_n11045_;
   wire new_n11041_;
   wire new_n11040_;
   wire new_n11039_;
   wire new_n11038_;
   wire new_n11037_;
   wire new_n11036_;
   wire new_n11035_;
   wire new_n11034_;
   wire new_n11027_;
   wire new_n11019_;
   wire new_n11018_;
   wire new_n11017_;
   wire new_n11015_;
   wire new_n11006_;
   wire new_n11005_;
   wire new_n11004_;
   wire new_n11003_;
   wire new_n11002_;
   wire new_n11001_;
   wire new_n11000_;
   wire new_n10999_;
   wire new_n10998_;
   wire new_n10997_;
   wire new_n10994_;
   wire new_n10993_;
   wire new_n10986_;
   wire new_n10985_;
   wire new_n10982_;
   wire new_n10981_;
   wire new_n10979_;
   wire new_n10978_;
   wire new_n10977_;
   wire new_n10976_;
   wire new_n10975_;
   wire new_n10974_;
   wire new_n10973_;
   wire new_n10972_;
   wire new_n10971_;
   wire new_n10969_;
   wire new_n10968_;
   wire new_n10963_;
   wire new_n10962_;
   wire new_n10955_;
   wire new_n10954_;
   wire new_n10952_;
   wire new_n10951_;
   wire new_n10950_;
   wire new_n10949_;
   wire new_n10948_;
   wire new_n10947_;
   wire new_n10946_;
   wire new_n10945_;
   wire new_n10944_;
   wire new_n10940_;
   wire new_n10939_;
   wire new_n10933_;
   wire new_n10932_;
   wire new_n10930_;
   wire new_n10929_;
   wire new_n10926_;
   wire new_n10925_;
   wire new_n10918_;
   wire new_n10917_;
   wire new_n10914_;
   wire new_n10913_;
   wire new_n10912_;
   wire new_n10911_;
   wire new_n10910_;
   wire new_n10909_;
   wire new_n10908_;
   wire new_n10907_;
   wire new_n10906_;
   wire new_n10903_;
   wire new_n10902_;
   wire new_n10896_;
   wire new_n10895_;
   wire new_n10893_;
   wire new_n10892_;
   wire new_n10890_;
   wire new_n10880_;
   wire new_n10879_;
   wire new_n10875_;
   wire new_n10874_;
   wire new_n10871_;
   wire new_n10869_;
   wire new_n10868_;
   wire new_n10867_;
   wire new_n10866_;
   wire new_n10865_;
   wire new_n10864_;
   wire new_n10863_;
   wire new_n10862_;
   wire new_n10861_;
   wire new_n10860_;
   wire new_n10857_;
   wire new_n10856_;
   wire new_n10855_;
   wire new_n10854_;
   wire new_n10853_;
   wire new_n10852_;
   wire new_n10851_;
   wire new_n10850_;
   wire new_n10849_;
   wire new_n10839_;
   wire new_n10838_;
   wire new_n10837_;
   wire new_n10836_;
   wire new_n10835_;
   wire new_n10834_;
   wire new_n10833_;
   wire new_n10832_;
   wire new_n10831_;
   wire new_n10830_;
   wire new_n10829_;
   wire new_n10828_;
   wire new_n10827_;
   wire new_n10826_;
   wire new_n10825_;
   wire new_n10824_;
   wire new_n10823_;
   wire new_n10822_;
   wire new_n10821_;
   wire new_n10820_;
   wire new_n10819_;
   wire new_n10818_;
   wire new_n10817_;
   wire new_n10816_;
   wire new_n10815_;
   wire new_n10811_;
   wire new_n10810_;
   wire new_n10805_;
   wire new_n10804_;
   wire new_n10803_;
   wire new_n10802_;
   wire new_n10801_;
   wire new_n10800_;
   wire new_n10799_;
   wire new_n10798_;
   wire new_n10797_;
   wire new_n10796_;
   wire new_n10795_;
   wire new_n10794_;
   wire new_n10793_;
   wire new_n10792_;
   wire new_n10785_;
   wire new_n10784_;
   wire new_n10783_;
   wire new_n10782_;
   wire new_n10781_;
   wire new_n10780_;
   wire new_n10779_;
   wire new_n10778_;
   wire new_n10777_;
   wire new_n10776_;
   wire new_n10775_;
   wire new_n10774_;
   wire new_n10767_;
   wire new_n10766_;
   wire new_n10765_;
   wire new_n10764_;
   wire new_n10761_;
   wire new_n10756_;
   wire new_n10755_;
   wire new_n10754_;
   wire new_n10753_;
   wire new_n10752_;
   wire new_n10751_;
   wire new_n10749_;
   wire new_n10748_;
   wire new_n10746_;
   wire new_n10745_;
   wire new_n10744_;
   wire new_n10743_;
   wire new_n10742_;
   wire new_n10741_;
   wire new_n10740_;
   wire new_n10739_;
   wire new_n10738_;
   wire new_n10737_;
   wire new_n10736_;
   wire new_n10735_;
   wire new_n10734_;
   wire new_n10733_;
   wire new_n10732_;
   wire new_n10730_;
   wire new_n10729_;
   wire new_n10726_;
   wire new_n10725_;
   wire new_n10721_;
   wire new_n10720_;
   wire new_n10712_;
   wire new_n10711_;
   wire new_n10707_;
   wire new_n10706_;
   wire new_n10704_;
   wire new_n10703_;
   wire new_n10702_;
   wire new_n10701_;
   wire new_n10692_;
   wire new_n10691_;
   wire new_n10690_;
   wire new_n10680_;
   wire new_n10679_;
   wire new_n10677_;
   wire new_n10673_;
   wire new_n10672_;
   wire new_n10666_;
   wire new_n10665_;
   wire new_n10660_;
   wire new_n10659_;
   wire new_n10658_;
   wire new_n10657_;
   wire new_n10656_;
   wire new_n10655_;
   wire new_n10654_;
   wire new_n10653_;
   wire new_n10652_;
   wire new_n10651_;
   wire new_n10650_;
   wire new_n10649_;
   wire new_n10648_;
   wire new_n10647_;
   wire new_n10642_;
   wire new_n10641_;
   wire new_n10640_;
   wire new_n10637_;
   wire new_n10636_;
   wire new_n10631_;
   wire new_n10628_;
   wire new_n10627_;
   wire new_n10626_;
   wire new_n10625_;
   wire new_n10624_;
   wire new_n10623_;
   wire new_n10622_;
   wire new_n10621_;
   wire new_n10620_;
   wire new_n10619_;
   wire new_n10618_;
   wire new_n10617_;
   wire new_n10616_;
   wire new_n10615_;
   wire new_n10608_;
   wire new_n10607_;
   wire new_n10606_;
   wire new_n10605_;
   wire new_n10600_;
   wire new_n10599_;
   wire new_n10598_;
   wire new_n10597_;
   wire new_n10595_;
   wire new_n10594_;
   wire new_n10593_;
   wire new_n10592_;
   wire new_n10591_;
   wire new_n10590_;
   wire new_n10589_;
   wire new_n10588_;
   wire new_n10587_;
   wire new_n10586_;
   wire new_n10585_;
   wire new_n10584_;
   wire new_n10583_;
   wire new_n10582_;
   wire new_n10579_;
   wire new_n10576_;
   wire new_n10575_;
   wire new_n10573_;
   wire new_n10572_;
   wire new_n10567_;
   wire new_n10566_;
   wire new_n10564_;
   wire new_n10559_;
   wire new_n10558_;
   wire new_n10557_;
   wire new_n10556_;
   wire new_n10555_;
   wire new_n10552_;
   wire new_n10551_;
   wire new_n10550_;
   wire new_n10549_;
   wire new_n10548_;
   wire new_n10547_;
   wire new_n10546_;
   wire new_n10545_;
   wire new_n10544_;
   wire new_n10543_;
   wire new_n10542_;
   wire new_n10541_;
   wire new_n10540_;
   wire new_n10539_;
   wire new_n10536_;
   wire new_n10535_;
   wire new_n10530_;
   wire new_n10529_;
   wire new_n10528_;
   wire new_n10527_;
   wire new_n10526_;
   wire new_n10525_;
   wire new_n10524_;
   wire new_n10522_;
   wire new_n10521_;
   wire new_n10517_;
   wire new_n10516_;
   wire new_n10515_;
   wire new_n10514_;
   wire new_n10506_;
   wire new_n10505_;
   wire new_n10499_;
   wire new_n10498_;
   wire new_n10497_;
   wire new_n10496_;
   wire new_n10495_;
   wire new_n10494_;
   wire new_n10493_;
   wire new_n10492_;
   wire new_n10491_;
   wire new_n10490_;
   wire new_n10489_;
   wire new_n10488_;
   wire new_n10487_;
   wire new_n10486_;
   wire new_n10479_;
   wire new_n10478_;
   wire new_n10476_;
   wire new_n10475_;
   wire new_n10473_;
   wire new_n10472_;
   wire new_n10469_;
   wire new_n10468_;
   wire new_n10464_;
   wire new_n10463_;
   wire new_n10460_;
   wire new_n10459_;
   wire new_n10458_;
   wire new_n10457_;
   wire new_n10456_;
   wire new_n10455_;
   wire new_n10454_;
   wire new_n10453_;
   wire new_n10452_;
   wire new_n10448_;
   wire new_n10447_;
   wire new_n10444_;
   wire new_n10443_;
   wire new_n10442_;
   wire new_n10441_;
   wire new_n10440_;
   wire new_n10439_;
   wire new_n10438_;
   wire new_n10437_;
   wire new_n10436_;
   wire new_n10428_;
   wire new_n10427_;
   wire new_n10425_;
   wire new_n10424_;
   wire new_n10422_;
   wire new_n10421_;
   wire new_n10419_;
   wire new_n10418_;
   wire new_n10417_;
   wire new_n10414_;
   wire new_n10413_;
   wire new_n10395_;
   wire new_n10394_;
   wire new_n10390_;
   wire new_n10389_;
   wire new_n10380_;
   wire new_n10379_;
   wire new_n10377_;
   wire new_n10376_;
   wire new_n10371_;
   wire new_n10368_;
   wire new_n10367_;
   wire new_n10364_;
   wire new_n10359_;
   wire new_n10354_;
   wire new_n10353_;
   wire new_n10352_;
   wire new_n10351_;
   wire new_n10350_;
   wire new_n10349_;
   wire new_n10348_;
   wire new_n10347_;
   wire new_n10346_;
   wire new_n10340_;
   wire new_n10339_;
   wire new_n10337_;
   wire new_n10336_;
   wire new_n10335_;
   wire new_n10325_;
   wire new_n10322_;
   wire new_n10314_;
   wire new_n10305_;
   wire new_n10303_;
   wire new_n10302_;
   wire new_n10301_;
   wire new_n10300_;
   wire new_n10299_;
   wire new_n10298_;
   wire new_n10297_;
   wire new_n10296_;
   wire new_n10295_;
   wire new_n10294_;
   wire new_n10293_;
   wire new_n10292_;
   wire new_n10291_;
   wire new_n10290_;
   wire new_n10284_;
   wire new_n10283_;
   wire new_n10281_;
   wire new_n10280_;
   wire new_n10279_;
   wire new_n10278_;
   wire new_n10277_;
   wire new_n10276_;
   wire new_n10275_;
   wire new_n10274_;
   wire new_n10273_;
   wire new_n10266_;
   wire new_n10265_;
   wire new_n10263_;
   wire new_n10262_;
   wire new_n10253_;
   wire new_n10252_;
   wire new_n10250_;
   wire new_n10249_;
   wire new_n10248_;
   wire new_n10247_;
   wire new_n10246_;
   wire new_n10245_;
   wire new_n10244_;
   wire new_n10242_;
   wire new_n10241_;
   wire new_n10240_;
   wire new_n10239_;
   wire new_n10238_;
   wire new_n10237_;
   wire new_n10234_;
   wire new_n10233_;
   wire new_n10232_;
   wire new_n10231_;
   wire new_n10230_;
   wire new_n10229_;
   wire new_n10228_;
   wire new_n10227_;
   wire new_n10226_;
   wire new_n10225_;
   wire new_n10222_;
   wire new_n10221_;
   wire new_n10216_;
   wire new_n10215_;
   wire new_n10198_;
   wire new_n10197_;
   wire new_n10193_;
   wire new_n10192_;
   wire new_n10189_;
   wire new_n10188_;
   wire new_n10185_;
   wire new_n10184_;
   wire new_n10183_;
   wire new_n10182_;
   wire new_n10181_;
   wire new_n10180_;
   wire new_n10179_;
   wire new_n10178_;
   wire new_n10177_;
   wire new_n10176_;
   wire new_n10175_;
   wire new_n10174_;
   wire new_n10173_;
   wire new_n10172_;
   wire new_n10163_;
   wire new_n10162_;
   wire new_n10159_;
   wire new_n10158_1_;
   wire new_n10157_;
   wire new_n10151_;
   wire new_n10150_1_;
   wire new_n10148_;
   wire new_n10147_;
   wire new_n10144_;
   wire new_n10143_;
   wire new_n10136_;
   wire new_n10135_;
   wire new_n10133_;
   wire new_n10132_1_;
   wire new_n10131_;
   wire new_n10130_;
   wire new_n10129_;
   wire new_n10126_;
   wire new_n10125_;
   wire new_n10121_;
   wire new_n10115_;
   wire new_n10114_;
   wire new_n10112_1_;
   wire new_n10111_;
   wire new_n10110_;
   wire new_n10106_;
   wire new_n10105_;
   wire new_n10104_;
   wire new_n10103_1_;
   wire new_n10102_;
   wire new_n10101_;
   wire new_n10100_;
   wire new_n10099_1_;
   wire new_n10098_;
   wire new_n10097_;
   wire new_n10095_;
   wire new_n10094_1_;
   wire new_n10093_;
   wire new_n10092_;
   wire new_n10091_;
   wire new_n10090_;
   wire new_n10089_1_;
   wire new_n10086_;
   wire new_n10085_;
   wire new_n10084_1_;
   wire new_n10076_;
   wire new_n10075_;
   wire new_n10068_;
   wire new_n10067_;
   wire new_n10064_;
   wire new_n10063_;
   wire new_n10058_;
   wire new_n10056_1_;
   wire new_n10055_;
   wire new_n10054_;
   wire new_n10053_;
   wire new_n10052_1_;
   wire new_n10051_;
   wire new_n10049_;
   wire new_n10047_1_;
   wire new_n10046_;
   wire new_n10045_;
   wire new_n10044_;
   wire new_n10043_;
   wire new_n10042_1_;
   wire new_n10041_;
   wire new_n10040_;
   wire new_n10039_;
   wire new_n10038_;
   wire new_n10035_;
   wire new_n10034_;
   wire new_n10031_;
   wire new_n10030_;
   wire new_n10028_1_;
   wire new_n10027_;
   wire new_n10025_;
   wire new_n10021_;
   wire new_n10010_1_;
   wire new_n10009_;
   wire new_n10008_;
   wire new_n10006_1_;
   wire new_n10005_;
   wire net_7807;
   wire net_7802;
   wire net_7799;
   wire net_7792;
   wire net_7790;
   wire net_7780;
   wire net_7779;
   wire net_7778;
   wire net_7777;
   wire net_7776;
   wire net_7775;
   wire net_7774;
   wire net_7773;
   wire net_7772;
   wire net_7771;
   wire net_7770;
   wire net_7769;
   wire net_7767;
   wire net_7766;
   wire net_7764;
   wire net_7762;
   wire net_7760;
   wire net_7758;
   wire net_7756;
   wire net_7754;
   wire net_7752;
   wire net_7750;
   wire net_7744;
   wire net_7743;
   wire net_7742;
   wire net_7741;
   wire net_7740;
   wire net_7739;
   wire net_7738;
   wire net_7737;
   wire net_7715;
   wire net_7714;
   wire net_7713;
   wire net_7712;
   wire net_7711;
   wire net_7710;
   wire net_7709;
   wire net_7708;
   wire net_7691;
   wire net_7680;
   wire net_7679;
   wire net_7678;
   wire net_7677;
   wire net_7676;
   wire net_7675;
   wire net_7674;
   wire net_7673;
   wire net_7672;
   wire net_7671;
   wire net_7670;
   wire net_7669;
   wire net_7668;
   wire net_7647;
   wire net_7646;
   wire net_7645;
   wire net_7644;
   wire net_7643;
   wire net_7642;
   wire net_7641;
   wire net_7640;
   wire net_7639;
   wire net_7638;
   wire net_7637;
   wire net_7636;
   wire net_7615;
   wire net_7614;
   wire net_7613;
   wire net_7612;
   wire net_7611;
   wire net_7610;
   wire net_7609;
   wire net_7608;
   wire net_7607;
   wire net_7606;
   wire net_7605;
   wire net_7604;
   wire net_7551;
   wire net_7550;
   wire net_7549;
   wire net_7548;
   wire net_7547;
   wire net_7546;
   wire net_7545;
   wire net_7544;
   wire net_7543;
   wire net_7542;
   wire net_7541;
   wire net_7540;
   wire net_7539;
   wire net_7538;
   wire net_7537;
   wire net_7536;
   wire net_7529;
   wire net_7528;
   wire net_7527;
   wire net_7526;
   wire net_7525;
   wire net_7524;
   wire net_7523;
   wire net_7522;
   wire net_7521;
   wire net_7520;
   wire net_7519;
   wire net_7518;
   wire net_7517;
   wire net_7496;
   wire net_7495;
   wire net_7494;
   wire net_7493;
   wire net_7492;
   wire net_7491;
   wire net_7490;
   wire net_7489;
   wire net_7488;
   wire net_7487;
   wire net_7486;
   wire net_7485;
   wire net_7464;
   wire net_7463;
   wire net_7462;
   wire net_7461;
   wire net_7460;
   wire net_7459;
   wire net_7458;
   wire net_7457;
   wire net_7456;
   wire net_7455;
   wire net_7454;
   wire net_7453;
   wire net_7400;
   wire net_7399;
   wire net_7398;
   wire net_7397;
   wire net_7396;
   wire net_7395;
   wire net_7394;
   wire net_7393;
   wire net_7392;
   wire net_7391;
   wire net_7390;
   wire net_7389;
   wire net_7388;
   wire net_7387;
   wire net_7386;
   wire net_7385;
   wire net_7378;
   wire net_7377;
   wire net_7376;
   wire net_7375;
   wire net_7374;
   wire net_7373;
   wire net_7372;
   wire net_7371;
   wire net_7370;
   wire net_7369;
   wire net_7368;
   wire net_7367;
   wire net_7366;
   wire net_7345;
   wire net_7344;
   wire net_7343;
   wire net_7342;
   wire net_7341;
   wire net_7340;
   wire net_7339;
   wire net_7338;
   wire net_7337;
   wire net_7336;
   wire net_7335;
   wire net_7334;
   wire net_7313;
   wire net_7312;
   wire net_7311;
   wire net_7310;
   wire net_7309;
   wire net_7308;
   wire net_7307;
   wire net_7306;
   wire net_7305;
   wire net_7304;
   wire net_7303;
   wire net_7302;
   wire net_7249;
   wire net_7248;
   wire net_7247;
   wire net_7246;
   wire net_7245;
   wire net_7244;
   wire net_7243;
   wire net_7242;
   wire net_7241;
   wire net_7240;
   wire net_7239;
   wire net_7238;
   wire net_7237;
   wire net_7236;
   wire net_7235;
   wire net_7234;
   wire net_7231;
   wire net_7226;
   wire net_7225;
   wire net_7224;
   wire net_7223;
   wire net_7222;
   wire net_7221;
   wire net_7220;
   wire net_7219;
   wire net_7218;
   wire net_7217;
   wire net_7216;
   wire net_7215;
   wire net_7214;
   wire net_7213;
   wire net_7212;
   wire net_7211;
   wire net_7210;
   wire net_7209;
   wire net_7208;
   wire net_7207;
   wire net_7206;
   wire net_7205;
   wire net_7204;
   wire net_7203;
   wire net_7202;
   wire net_7201;
   wire net_7200;
   wire net_7199;
   wire net_7198;
   wire net_7197;
   wire net_7196;
   wire net_7195;
   wire net_7194;
   wire net_7193;
   wire net_7192;
   wire net_7191;
   wire net_7190;
   wire net_7189;
   wire net_7188;
   wire net_7187;
   wire net_7186;
   wire net_7185;
   wire net_7184;
   wire net_7183;
   wire net_7182;
   wire net_7181;
   wire net_7180;
   wire net_7179;
   wire net_7178;
   wire net_7177;
   wire net_7176;
   wire net_7175;
   wire net_7174;
   wire net_7173;
   wire net_7172;
   wire net_7171;
   wire net_7170;
   wire net_7169;
   wire net_7168;
   wire net_7167;
   wire net_7166;
   wire net_7165;
   wire net_7164;
   wire net_7163;
   wire net_7162;
   wire net_7161;
   wire net_7160;
   wire net_7159;
   wire net_7158;
   wire net_7157;
   wire net_7156;
   wire net_7155;
   wire net_7154;
   wire net_7153;
   wire net_7152;
   wire net_7151;
   wire net_7150;
   wire net_7149;
   wire net_7148;
   wire net_7147;
   wire net_7146;
   wire net_7145;
   wire net_7144;
   wire net_7143;
   wire net_7142;
   wire net_7141;
   wire net_7140;
   wire net_7139;
   wire net_7138;
   wire net_7137;
   wire net_7136;
   wire net_7135;
   wire net_7134;
   wire net_7133;
   wire net_7132;
   wire net_7131;
   wire net_7130;
   wire net_7129;
   wire net_7128;
   wire net_7127;
   wire net_7126;
   wire net_7125;
   wire net_7124;
   wire net_7123;
   wire net_7122;
   wire net_7121;
   wire net_7120;
   wire net_7119;
   wire net_7118;
   wire net_7117;
   wire net_7116;
   wire net_7115;
   wire net_7114;
   wire net_7113;
   wire net_7112;
   wire net_7111;
   wire net_7110;
   wire net_7109;
   wire net_7108;
   wire net_7107;
   wire net_7106;
   wire net_7105;
   wire net_7104;
   wire net_7103;
   wire net_7102;
   wire net_7101;
   wire net_7100;
   wire net_7099;
   wire net_7096;
   wire net_7091;
   wire net_7090;
   wire net_7089;
   wire net_7088;
   wire net_7087;
   wire net_7086;
   wire net_7085;
   wire net_7084;
   wire net_7083;
   wire net_7082;
   wire net_7081;
   wire net_7080;
   wire net_7079;
   wire net_7078;
   wire net_7077;
   wire net_7076;
   wire net_7075;
   wire net_7074;
   wire net_7073;
   wire net_7072;
   wire net_7071;
   wire net_7070;
   wire net_7069;
   wire net_7068;
   wire net_7067;
   wire net_7066;
   wire net_7065;
   wire net_7064;
   wire net_7063;
   wire net_7062;
   wire net_7061;
   wire net_7060;
   wire net_7059;
   wire net_7058;
   wire net_7057;
   wire net_7056;
   wire net_7055;
   wire net_7054;
   wire net_7053;
   wire net_7052;
   wire net_7051;
   wire net_7050;
   wire net_7049;
   wire net_7048;
   wire net_7047;
   wire net_7046;
   wire net_7045;
   wire net_7044;
   wire net_7043;
   wire net_7042;
   wire net_7041;
   wire net_7040;
   wire net_7039;
   wire net_7038;
   wire net_7037;
   wire net_7036;
   wire net_7035;
   wire net_7034;
   wire net_7033;
   wire net_7032;
   wire net_7031;
   wire net_7030;
   wire net_7029;
   wire net_7028;
   wire net_7027;
   wire net_7026;
   wire net_7025;
   wire net_7024;
   wire net_7023;
   wire net_7022;
   wire net_7021;
   wire net_7020;
   wire net_7019;
   wire net_7018;
   wire net_7017;
   wire net_7016;
   wire net_7015;
   wire net_7014;
   wire net_7013;
   wire net_7012;
   wire net_7011;
   wire net_7010;
   wire net_7009;
   wire net_7008;
   wire net_7007;
   wire net_7006;
   wire net_7005;
   wire net_7004;
   wire net_7003;
   wire net_7002;
   wire net_7001;
   wire net_7000;
   wire net_6999;
   wire net_6998;
   wire net_6997;
   wire net_6996;
   wire net_6995;
   wire net_6994;
   wire net_6993;
   wire net_6992;
   wire net_6991;
   wire net_6990;
   wire net_6989;
   wire net_6988;
   wire net_6987;
   wire net_6986;
   wire net_6985;
   wire net_6984;
   wire net_6983;
   wire net_6982;
   wire net_6981;
   wire net_6980;
   wire net_6979;
   wire net_6978;
   wire net_6977;
   wire net_6976;
   wire net_6975;
   wire net_6974;
   wire net_6973;
   wire net_6972;
   wire net_6971;
   wire net_6970;
   wire net_6969;
   wire net_6968;
   wire net_6967;
   wire net_6966;
   wire net_6965;
   wire net_6964;
   wire net_6961;
   wire net_6956;
   wire net_6955;
   wire net_6954;
   wire net_6953;
   wire net_6952;
   wire net_6951;
   wire net_6950;
   wire net_6949;
   wire net_6948;
   wire net_6947;
   wire net_6946;
   wire net_6945;
   wire net_6944;
   wire net_6943;
   wire net_6942;
   wire net_6941;
   wire net_6940;
   wire net_6939;
   wire net_6938;
   wire net_6937;
   wire net_6936;
   wire net_6935;
   wire net_6934;
   wire net_6933;
   wire net_6932;
   wire net_6931;
   wire net_6930;
   wire net_6929;
   wire net_6928;
   wire net_6927;
   wire net_6926;
   wire net_6925;
   wire net_6924;
   wire net_6923;
   wire net_6922;
   wire net_6921;
   wire net_6920;
   wire net_6919;
   wire net_6918;
   wire net_6917;
   wire net_6916;
   wire net_6915;
   wire net_6914;
   wire net_6913;
   wire net_6912;
   wire net_6911;
   wire net_6910;
   wire net_6909;
   wire net_6908;
   wire net_6907;
   wire net_6906;
   wire net_6905;
   wire net_6904;
   wire net_6903;
   wire net_6902;
   wire net_6901;
   wire net_6900;
   wire net_6899;
   wire net_6898;
   wire net_6897;
   wire net_6896;
   wire net_6895;
   wire net_6894;
   wire net_6893;
   wire net_6892;
   wire net_6891;
   wire net_6890;
   wire net_6889;
   wire net_6888;
   wire net_6887;
   wire net_6886;
   wire net_6885;
   wire net_6884;
   wire net_6883;
   wire net_6882;
   wire net_6881;
   wire net_6880;
   wire net_6879;
   wire net_6878;
   wire net_6877;
   wire net_6876;
   wire net_6875;
   wire net_6874;
   wire net_6873;
   wire net_6872;
   wire net_6871;
   wire net_6870;
   wire net_6869;
   wire net_6868;
   wire net_6867;
   wire net_6866;
   wire net_6865;
   wire net_6864;
   wire net_6863;
   wire net_6862;
   wire net_6861;
   wire net_6860;
   wire net_6859;
   wire net_6858;
   wire net_6857;
   wire net_6856;
   wire net_6855;
   wire net_6854;
   wire net_6853;
   wire net_6852;
   wire net_6851;
   wire net_6850;
   wire net_6849;
   wire net_6848;
   wire net_6847;
   wire net_6846;
   wire net_6845;
   wire net_6844;
   wire net_6843;
   wire net_6842;
   wire net_6841;
   wire net_6840;
   wire net_6839;
   wire net_6838;
   wire net_6837;
   wire net_6836;
   wire net_6835;
   wire net_6834;
   wire net_6833;
   wire net_6832;
   wire net_6831;
   wire net_6830;
   wire net_6829;
   wire net_6826;
   wire net_6821;
   wire net_6820;
   wire net_6819;
   wire net_6818;
   wire net_6817;
   wire net_6816;
   wire net_6815;
   wire net_6814;
   wire net_6813;
   wire net_6812;
   wire net_6811;
   wire net_6810;
   wire net_6809;
   wire net_6808;
   wire net_6807;
   wire net_6806;
   wire net_6805;
   wire net_6804;
   wire net_6803;
   wire net_6802;
   wire net_6801;
   wire net_6800;
   wire net_6799;
   wire net_6798;
   wire net_6797;
   wire net_6796;
   wire net_6795;
   wire net_6794;
   wire net_6793;
   wire net_6792;
   wire net_6791;
   wire net_6790;
   wire net_6789;
   wire net_6788;
   wire net_6787;
   wire net_6786;
   wire net_6785;
   wire net_6784;
   wire net_6783;
   wire net_6782;
   wire net_6781;
   wire net_6780;
   wire net_6779;
   wire net_6778;
   wire net_6777;
   wire net_6776;
   wire net_6775;
   wire net_6774;
   wire net_6773;
   wire net_6772;
   wire net_6771;
   wire net_6770;
   wire net_6769;
   wire net_6768;
   wire net_6767;
   wire net_6766;
   wire net_6765;
   wire net_6764;
   wire net_6763;
   wire net_6762;
   wire net_6761;
   wire net_6760;
   wire net_6759;
   wire net_6758;
   wire net_6757;
   wire net_6756;
   wire net_6755;
   wire net_6754;
   wire net_6753;
   wire net_6752;
   wire net_6751;
   wire net_6750;
   wire net_6749;
   wire net_6748;
   wire net_6747;
   wire net_6746;
   wire net_6745;
   wire net_6744;
   wire net_6743;
   wire net_6742;
   wire net_6741;
   wire net_6740;
   wire net_6739;
   wire net_6738;
   wire net_6737;
   wire net_6736;
   wire net_6735;
   wire net_6734;
   wire net_6733;
   wire net_6732;
   wire net_6731;
   wire net_6730;
   wire net_6729;
   wire net_6728;
   wire net_6727;
   wire net_6726;
   wire net_6725;
   wire net_6724;
   wire net_6723;
   wire net_6722;
   wire net_6721;
   wire net_6720;
   wire net_6719;
   wire net_6718;
   wire net_6717;
   wire net_6716;
   wire net_6715;
   wire net_6714;
   wire net_6713;
   wire net_6712;
   wire net_6711;
   wire net_6710;
   wire net_6709;
   wire net_6708;
   wire net_6707;
   wire net_6706;
   wire net_6705;
   wire net_6704;
   wire net_6703;
   wire net_6702;
   wire net_6701;
   wire net_6700;
   wire net_6699;
   wire net_6698;
   wire net_6697;
   wire net_6696;
   wire net_6695;
   wire net_6694;
   wire net_6691;
   wire net_6686;
   wire net_6685;
   wire net_6684;
   wire net_6683;
   wire net_6682;
   wire net_6681;
   wire net_6680;
   wire net_6679;
   wire net_6678;
   wire net_6677;
   wire net_6676;
   wire net_6675;
   wire net_6674;
   wire net_6673;
   wire net_6672;
   wire net_6671;
   wire net_6670;
   wire net_6669;
   wire net_6668;
   wire net_6667;
   wire net_6666;
   wire net_6665;
   wire net_6664;
   wire net_6663;
   wire net_6662;
   wire net_6661;
   wire net_6660;
   wire net_6659;
   wire net_6658;
   wire net_6657;
   wire net_6656;
   wire net_6655;
   wire net_6654;
   wire net_6653;
   wire net_6652;
   wire net_6651;
   wire net_6650;
   wire net_6649;
   wire net_6648;
   wire net_6647;
   wire net_6646;
   wire net_6645;
   wire net_6644;
   wire net_6643;
   wire net_6642;
   wire net_6641;
   wire net_6640;
   wire net_6639;
   wire net_6638;
   wire net_6637;
   wire net_6636;
   wire net_6635;
   wire net_6634;
   wire net_6633;
   wire net_6632;
   wire net_6631;
   wire net_6630;
   wire net_6629;
   wire net_6628;
   wire net_6627;
   wire net_6626;
   wire net_6625;
   wire net_6624;
   wire net_6623;
   wire net_6622;
   wire net_6621;
   wire net_6620;
   wire net_6619;
   wire net_6618;
   wire net_6617;
   wire net_6616;
   wire net_6615;
   wire net_6614;
   wire net_6613;
   wire net_6612;
   wire net_6611;
   wire net_6610;
   wire net_6609;
   wire net_6608;
   wire net_6607;
   wire net_6606;
   wire net_6605;
   wire net_6604;
   wire net_6603;
   wire net_6602;
   wire net_6601;
   wire net_6600;
   wire net_6599;
   wire net_6598;
   wire net_6597;
   wire net_6596;
   wire net_6595;
   wire net_6594;
   wire net_6593;
   wire net_6592;
   wire net_6591;
   wire net_6590;
   wire net_6589;
   wire net_6588;
   wire net_6587;
   wire net_6586;
   wire net_6585;
   wire net_6584;
   wire net_6583;
   wire net_6582;
   wire net_6581;
   wire net_6580;
   wire net_6579;
   wire net_6578;
   wire net_6577;
   wire net_6576;
   wire net_6575;
   wire net_6574;
   wire net_6573;
   wire net_6572;
   wire net_6571;
   wire net_6570;
   wire net_6569;
   wire net_6568;
   wire net_6567;
   wire net_6566;
   wire net_6565;
   wire net_6564;
   wire net_6563;
   wire net_6562;
   wire net_6561;
   wire net_6560;
   wire net_6559;
   wire net_6556;
   wire net_6551;
   wire net_6550;
   wire net_6549;
   wire net_6548;
   wire net_6547;
   wire net_6546;
   wire net_6545;
   wire net_6544;
   wire net_6543;
   wire net_6542;
   wire net_6541;
   wire net_6540;
   wire net_6539;
   wire net_6538;
   wire net_6537;
   wire net_6536;
   wire net_6535;
   wire net_6534;
   wire net_6533;
   wire net_6532;
   wire net_6531;
   wire net_6530;
   wire net_6529;
   wire net_6528;
   wire net_6527;
   wire net_6526;
   wire net_6525;
   wire net_6524;
   wire net_6523;
   wire net_6522;
   wire net_6521;
   wire net_6520;
   wire net_6519;
   wire net_6518;
   wire net_6517;
   wire net_6516;
   wire net_6515;
   wire net_6514;
   wire net_6513;
   wire net_6512;
   wire net_6511;
   wire net_6510;
   wire net_6509;
   wire net_6508;
   wire net_6507;
   wire net_6506;
   wire net_6505;
   wire net_6504;
   wire net_6503;
   wire net_6502;
   wire net_6501;
   wire net_6500;
   wire net_6499;
   wire net_6498;
   wire net_6497;
   wire net_6496;
   wire net_6495;
   wire net_6494;
   wire net_6493;
   wire net_6492;
   wire net_6491;
   wire net_6490;
   wire net_6489;
   wire net_6488;
   wire net_6487;
   wire net_6486;
   wire net_6485;
   wire net_6484;
   wire net_6483;
   wire net_6482;
   wire net_6481;
   wire net_6480;
   wire net_6479;
   wire net_6478;
   wire net_6477;
   wire net_6476;
   wire net_6475;
   wire net_6474;
   wire net_6473;
   wire net_6472;
   wire net_6471;
   wire net_6470;
   wire net_6469;
   wire net_6468;
   wire net_6467;
   wire net_6466;
   wire net_6465;
   wire net_6464;
   wire net_6463;
   wire net_6462;
   wire net_6461;
   wire net_6460;
   wire net_6459;
   wire net_6458;
   wire net_6457;
   wire net_6456;
   wire net_6455;
   wire net_6454;
   wire net_6453;
   wire net_6452;
   wire net_6451;
   wire net_6450;
   wire net_6449;
   wire net_6448;
   wire net_6447;
   wire net_6446;
   wire net_6445;
   wire net_6444;
   wire net_6443;
   wire net_6442;
   wire net_6441;
   wire net_6440;
   wire net_6439;
   wire net_6438;
   wire net_6437;
   wire net_6436;
   wire net_6435;
   wire net_6434;
   wire net_6433;
   wire net_6432;
   wire net_6431;
   wire net_6430;
   wire net_6429;
   wire net_6428;
   wire net_6427;
   wire net_6426;
   wire net_6425;
   wire net_6424;
   wire net_6417;
   wire net_6416;
   wire net_6412;
   wire net_6403;
   wire net_6400;
   wire net_6399;
   wire net_6398;
   wire net_6397;
   wire net_6396;
   wire net_6395;
   wire net_6394;
   wire net_6393;
   wire net_6392;
   wire net_6391;
   wire net_6390;
   wire net_6389;
   wire net_6388;
   wire net_6387;
   wire net_6386;
   wire net_6385;
   wire net_6384;
   wire net_6383;
   wire net_6382;
   wire net_6381;
   wire net_6380;
   wire net_6379;
   wire net_6378;
   wire net_6377;
   wire net_6376;
   wire net_6375;
   wire net_6374;
   wire net_6373;
   wire net_6372;
   wire net_6371;
   wire net_6370;
   wire net_6369;
   wire net_6368;
   wire net_6367;
   wire net_6366;
   wire net_6365;
   wire net_6364;
   wire net_6363;
   wire net_6362;
   wire net_6361;
   wire net_6360;
   wire net_6359;
   wire net_6358;
   wire net_6357;
   wire net_6356;
   wire net_6355;
   wire net_6354;
   wire net_6353;
   wire net_6352;
   wire net_6351;
   wire net_6350;
   wire net_6349;
   wire net_6348;
   wire net_6347;
   wire net_6346;
   wire net_6345;
   wire net_6344;
   wire net_6343;
   wire net_6342;
   wire net_6341;
   wire net_6340;
   wire net_6339;
   wire net_6338;
   wire net_6337;
   wire net_6336;
   wire net_6335;
   wire net_6334;
   wire net_6333;
   wire net_6332;
   wire net_6331;
   wire net_6330;
   wire net_6329;
   wire net_6328;
   wire net_6327;
   wire net_6326;
   wire net_6325;
   wire net_6324;
   wire net_6323;
   wire net_6322;
   wire net_6321;
   wire net_6320;
   wire net_6318;
   wire net_6317;
   wire net_6316;
   wire net_6315;
   wire net_6314;
   wire net_6313;
   wire net_6312;
   wire net_6311;
   wire net_6310;
   wire net_6309;
   wire net_6308;
   wire net_6307;
   wire net_6306;
   wire net_6305;
   wire net_6304;
   wire net_6303;
   wire net_6302;
   wire net_6301;
   wire net_6300;
   wire net_6299;
   wire net_6279;
   wire net_6278;
   wire net_6277;
   wire net_6276;
   wire net_6275;
   wire net_6274;
   wire net_6273;
   wire net_6272;
   wire net_6271;
   wire net_6270;
   wire net_6269;
   wire net_6268;
   wire net_6267;
   wire net_6266;
   wire net_6265;
   wire net_6264;
   wire net_6263;
   wire net_6262;
   wire net_6261;
   wire net_6260;
   wire net_6258;
   wire net_6257;
   wire net_6256;
   wire net_6255;
   wire net_6254;
   wire net_6253;
   wire net_6252;
   wire net_6251;
   wire net_6250;
   wire net_6249;
   wire net_6248;
   wire net_6247;
   wire net_6246;
   wire net_6245;
   wire net_6244;
   wire net_6243;
   wire net_6242;
   wire net_6241;
   wire net_6240;
   wire net_6238;
   wire net_6237;
   wire net_6236;
   wire net_6235;
   wire net_6234;
   wire net_6233;
   wire net_6232;
   wire net_6231;
   wire net_6230;
   wire net_6229;
   wire net_6228;
   wire net_6227;
   wire net_6226;
   wire net_6225;
   wire net_6224;
   wire net_6223;
   wire net_6218;
   wire net_6217;
   wire net_6216;
   wire net_6215;
   wire net_6214;
   wire net_6213;
   wire net_6212;
   wire net_6211;
   wire net_6198;
   wire net_6197;
   wire net_6196;
   wire net_6195;
   wire net_6193;
   wire net_6192;
   wire net_6191;
   wire net_6190;
   wire net_6061;
   wire net_6060;
   wire net_6059;
   wire net_6058;
   wire net_6057;
   wire net_6056;
   wire net_6055;
   wire net_6054;
   wire net_6053;
   wire net_6047;
   wire net_6046;
   wire net_6036;
   wire net_6035;
   wire net_6025;
   wire net_6024;
   wire net_6014;
   wire net_6013;
   wire net_6003;
   wire net_5992;
   wire net_5861;
   wire net_5860;
   wire net_5858;
   wire net_5849;
   wire net_391;
   wire net_390;
   wire net_389;
   wire net_388;
   wire net_387;
   wire net_386;
   wire net_385;
   wire net_384;
   wire net_383;
   wire net_382;
   wire net_381;
   wire net_380;
   wire net_379;
   wire net_378;
   wire net_377;
   wire net_376;
   wire net_375;
   wire net_374;
   wire net_373;
   wire net_372;
   wire net_371;
   wire net_370;
   wire net_369;
   wire net_368;
   wire net_367;
   wire net_366;
   wire net_365;
   wire net_364;
   wire net_363;
   wire net_362;
   wire net_361;
   wire net_360;
   wire net_359;
   wire net_358;
   wire net_357;
   wire net_356;
   wire net_355;
   wire net_354;
   wire net_353;
   wire net_352;
   wire net_351;
   wire net_350;
   wire net_349;
   wire net_348;
   wire net_347;
   wire net_346;
   wire net_345;
   wire net_344;
   wire net_343;
   wire net_342;
   wire net_341;
   wire net_340;
   wire net_339;
   wire net_338;
   wire net_337;
   wire net_336;
   wire net_335;
   wire net_334;
   wire net_333;
   wire net_332;
   wire net_331;
   wire net_330;
   wire net_329;
   wire net_328;
   wire net_327;
   wire net_326;
   wire net_325;
   wire net_324;
   wire net_323;
   wire net_322;
   wire net_321;
   wire net_320;
   wire net_319;
   wire net_318;
   wire net_317;
   wire net_316;
   wire net_315;
   wire net_314;
   wire net_313;
   wire net_312;
   wire net_311;
   wire net_310;
   wire net_309;
   wire net_308;
   wire net_307;
   wire net_306;
   wire net_305;
   wire net_304;
   wire net_303;
   wire net_302;
   wire net_301;
   wire net_300;
   wire net_297;
   wire net_296;
   wire net_286;
   wire net_285;
   wire net_275;
   wire net_274;
   wire net_261;
   wire net_260;
   wire net_259;
   wire net_258;
   wire net_257;
   wire net_256;
   wire net_255;
   wire net_254;
   wire net_253;
   wire net_252;
   wire net_251;
   wire net_250;
   wire net_249;
   wire net_248;
   wire net_247;
   wire net_246;
   wire net_245;
   wire net_244;
   wire net_243;
   wire net_242;
   wire net_241;
   wire net_240;
   wire net_239;
   wire net_238;
   wire net_237;
   wire net_236;
   wire net_235;
   wire net_234;
   wire net_233;
   wire net_232;
   wire net_231;
   wire net_230;
   wire net_224;
   wire net_223;
   wire net_222;
   wire net_220;
   wire net_219;
   wire net_218;
   wire net_216;
   wire net_208;
   wire net_207;
   wire net_206;
   wire net_205;
   wire net_204;
   wire net_203;
   wire net_202;
   wire net_200;
   wire net_199;
   wire net_198;
   wire net_197;
   wire net_196;
   wire net_195;
   wire net_194;
   wire net_187;
   wire net_186;
   wire net_185;
   wire net_183;
   wire net_182;
   wire net_181;
   wire net_179;
   wire net_171;
   wire net_170;
   wire net_169;
   wire net_168;
   wire net_167;
   wire net_166;
   wire net_165;
   wire net_164;
   wire net_163;
   wire net_162;
   wire net_161;
   wire net_160;
   wire net_159;
   wire net_158;
   wire net_157;
   wire net_156;
   wire net_155;
   wire net_153;
   wire net_152;
   wire net_151;
   wire net_150;
   wire net_149;
   wire net_148;
   wire net_147;
   wire net_146;
   wire net_145;
   wire net_144;
   wire net_143;
   wire net_142;
   wire net_141;
   wire net_140;
   wire net_139;
   wire net_138;
   wire net_137;
   wire net_136;
   wire net_135;
   wire net_134;
   wire net_133;
   wire net_132;
   wire net_131;
   wire net_130;
   wire n9997;
   wire n9992;
   wire n9988;
   wire n9985;
   wire n9981;
   wire n9976;
   wire n9971;
   wire n9966;
   wire n9961;
   wire n9957;
   wire n9953;
   wire n995;
   wire n9949;
   wire n9944;
   wire n9939;
   wire n9935;
   wire n9930;
   wire n9926;
   wire n9923;
   wire n9918;
   wire n9914;
   wire n9911;
   wire n9907;
   wire n9902;
   wire n990;
   wire n9899;
   wire n9894;
   wire n9889;
   wire n9885;
   wire n9880;
   wire n9875;
   wire n9871;
   wire n9867;
   wire n9863;
   wire n9858;
   wire n9853;
   wire n985;
   wire n9849;
   wire n9844;
   wire n9840;
   wire n9837;
   wire n9833;
   wire n9828;
   wire n9824;
   wire n9819;
   wire n9814;
   wire n981;
   wire n9809;
   wire n9805;
   wire n9801;
   wire n9796;
   wire n9792;
   wire n9787;
   wire n9783;
   wire n9778;
   wire n9773;
   wire n9768;
   wire n9763;
   wire n976;
   wire n9758;
   wire n9754;
   wire n9750;
   wire n9746;
   wire n9742;
   wire n9737;
   wire n9733;
   wire n9729;
   wire n9724;
   wire n9719;
   wire n9714;
   wire n971;
   wire n9709;
   wire n9704;
   wire n9700;
   wire n9695;
   wire n9692;
   wire n9687;
   wire n9683;
   wire n9678;
   wire n9673;
   wire n9668;
   wire n9664;
   wire n9660;
   wire n966;
   wire n9655;
   wire n9651;
   wire n9647;
   wire n9642;
   wire n9638;
   wire n9633;
   wire n9628;
   wire n9624;
   wire n9620;
   wire n9616;
   wire n9611;
   wire n961;
   wire n9606;
   wire n9602;
   wire n9597;
   wire n9592;
   wire n9588;
   wire n9583;
   wire n9579;
   wire n9574;
   wire n9569;
   wire n9564;
   wire n956;
   wire n9559;
   wire n9554;
   wire n9549;
   wire n9546;
   wire n9541;
   wire n9537;
   wire n9533;
   wire n953;
   wire n9528;
   wire n9525;
   wire n9520;
   wire n9517;
   wire n9512;
   wire n9507;
   wire n9502;
   wire n9497;
   wire n9492;
   wire n9487;
   wire n9483;
   wire n948;
   wire n9478;
   wire n9475;
   wire n9470;
   wire n9467;
   wire n9462;
   wire n9459;
   wire n9454;
   wire n9449;
   wire n9445;
   wire n9441;
   wire n944;
   wire n9436;
   wire n9431;
   wire n9428;
   wire n9425;
   wire n9420;
   wire n9415;
   wire n9410;
   wire n9405;
   wire n9402;
   wire n940;
   wire n9398;
   wire n9393;
   wire n9390;
   wire n9385;
   wire n9381;
   wire n9377;
   wire n9373;
   wire n9370;
   wire n9365;
   wire n9361;
   wire n9356;
   wire n9352;
   wire n935;
   wire n9348;
   wire n9343;
   wire n9339;
   wire n9335;
   wire n9330;
   wire n9326;
   wire n9321;
   wire n9316;
   wire n9312;
   wire n9307;
   wire n9302;
   wire n930;
   wire n9298;
   wire n9294;
   wire n9290;
   wire n9287;
   wire n9282;
   wire n9277;
   wire n9272;
   wire n9267;
   wire n9263;
   wire n9258;
   wire n9254;
   wire n9250;
   wire n925;
   wire n9245;
   wire n9242;
   wire n9238;
   wire n9233;
   wire n9228;
   wire n9225;
   wire n9220;
   wire n9215;
   wire n9211;
   wire n9206;
   wire n9201;
   wire n920;
   wire n9196;
   wire n9192;
   wire n9187;
   wire n9182;
   wire n9178;
   wire n9173;
   wire n9169;
   wire n9164;
   wire n9160;
   wire n916;
   wire n9156;
   wire n9151;
   wire n9146;
   wire n9143;
   wire n9138;
   wire n9134;
   wire n9129;
   wire n9124;
   wire n9120;
   wire n9115;
   wire n9110;
   wire n911;
   wire n9106;
   wire n9101;
   wire n9096;
   wire n9091;
   wire n9086;
   wire n9082;
   wire n9079;
   wire n9074;
   wire n907;
   wire n9069;
   wire n9065;
   wire n9060;
   wire n9057;
   wire n9052;
   wire n9047;
   wire n9042;
   wire n9037;
   wire n9034;
   wire n9030;
   wire n903;
   wire n9025;
   wire n9022;
   wire n9017;
   wire n9014;
   wire n9010;
   wire n9005;
   wire n9000;
   wire n8995;
   wire n8990;
   wire n899;
   wire n8986;
   wire n8981;
   wire n8976;
   wire n8971;
   wire n8967;
   wire n8963;
   wire n8958;
   wire n8953;
   wire n8948;
   wire n8943;
   wire n894;
   wire n8939;
   wire n8934;
   wire n8931;
   wire n8926;
   wire n8922;
   wire n8917;
   wire n8912;
   wire n8908;
   wire n8903;
   wire n890;
   wire n8899;
   wire n8895;
   wire n8891;
   wire n8886;
   wire n8882;
   wire n8877;
   wire n8873;
   wire n8869;
   wire n8864;
   wire n8860;
   wire n8855;
   wire n8850;
   wire n885;
   wire n8845;
   wire n8840;
   wire n8835;
   wire n8831;
   wire n8826;
   wire n8823;
   wire n8818;
   wire n8813;
   wire n8809;
   wire n8805;
   wire n8800;
   wire n880;
   wire n8797;
   wire n8793;
   wire n8788;
   wire n8784;
   wire n8780;
   wire n8775;
   wire n8771;
   wire n8767;
   wire n8762;
   wire n8757;
   wire n8753;
   wire n875;
   wire n8748;
   wire n8743;
   wire n8739;
   wire n8734;
   wire n8730;
   wire n8725;
   wire n8720;
   wire n8715;
   wire n8711;
   wire n8708;
   wire n8703;
   wire n870;
   wire n8698;
   wire n8694;
   wire n8689;
   wire n8685;
   wire n8681;
   wire n8676;
   wire n8671;
   wire n867;
   wire n8666;
   wire n8662;
   wire n8658;
   wire n8654;
   wire n8650;
   wire n8645;
   wire n8641;
   wire n8637;
   wire n8632;
   wire n8628;
   wire n8625;
   wire n8621;
   wire n862;
   wire n8616;
   wire n8612;
   wire n8607;
   wire n8602;
   wire n8598;
   wire n8593;
   wire n8588;
   wire n8583;
   wire n8578;
   wire n8575;
   wire n8570;
   wire n857;
   wire n8565;
   wire n8561;
   wire n8557;
   wire n8552;
   wire n8549;
   wire n8544;
   wire n8540;
   wire n854;
   wire n8535;
   wire n8531;
   wire n8526;
   wire n8522;
   wire n8517;
   wire n8513;
   wire n8508;
   wire n8504;
   wire n8499;
   wire n8494;
   wire n8491;
   wire n849;
   wire n8486;
   wire n8481;
   wire n8477;
   wire n8472;
   wire n8467;
   wire n8464;
   wire n8459;
   wire n8455;
   wire n8451;
   wire n8447;
   wire n8443;
   wire n844;
   wire n8438;
   wire n8435;
   wire n8430;
   wire n8426;
   wire n8422;
   wire n8418;
   wire n8415;
   wire n8410;
   wire n8405;
   wire n8401;
   wire n8396;
   wire n8392;
   wire n839;
   wire n8387;
   wire n8382;
   wire n8377;
   wire n8372;
   wire n8367;
   wire n8362;
   wire n8359;
   wire n8354;
   wire n8350;
   wire n8345;
   wire n8340;
   wire n834;
   wire n8337;
   wire n8334;
   wire n8329;
   wire n8324;
   wire n8320;
   wire n8316;
   wire n8311;
   wire n8307;
   wire n8303;
   wire n830;
   wire n8299;
   wire n8294;
   wire n8289;
   wire n8284;
   wire n8280;
   wire n8276;
   wire n8271;
   wire n8266;
   wire n8262;
   wire n8258;
   wire n8253;
   wire n825;
   wire n8249;
   wire n8245;
   wire n8241;
   wire n8237;
   wire n8232;
   wire n8228;
   wire n8224;
   wire n8220;
   wire n8216;
   wire n8211;
   wire n8206;
   wire n8202;
   wire n820;
   wire n8197;
   wire n8192;
   wire n8188;
   wire n8183;
   wire n8179;
   wire n8174;
   wire n8170;
   wire n8166;
   wire n8161;
   wire n8156;
   wire n8152;
   wire n815;
   wire n8147;
   wire n8144;
   wire n8140;
   wire n8135;
   wire n8130;
   wire n8125;
   wire n8121;
   wire n8116;
   wire n8112;
   wire n811;
   wire n8107;
   wire n8102;
   wire n8097;
   wire n8092;
   wire n8088;
   wire n8085;
   wire n8080;
   wire n8075;
   wire n8072;
   wire n8067;
   wire n8064;
   wire n806;
   wire n8059;
   wire n8056;
   wire n8051;
   wire n8047;
   wire n8042;
   wire n8038;
   wire n8033;
   wire n8028;
   wire n8024;
   wire n802;
   wire n8019;
   wire n8015;
   wire n8010;
   wire n8005;
   wire n8002;
   wire n7997;
   wire n7994;
   wire n7989;
   wire n7985;
   wire n7980;
   wire n798;
   wire n7975;
   wire n7970;
   wire n7967;
   wire n7962;
   wire n7958;
   wire n7955;
   wire n7950;
   wire n7945;
   wire n7942;
   wire n7937;
   wire n7933;
   wire n793;
   wire n7929;
   wire n7924;
   wire n7920;
   wire n7916;
   wire n7911;
   wire n7906;
   wire n7902;
   wire n7897;
   wire n7893;
   wire n7888;
   wire n7883;
   wire n788;
   wire n7878;
   wire n7875;
   wire n7871;
   wire n7867;
   wire n7863;
   wire n7858;
   wire n7853;
   wire n7848;
   wire n7845;
   wire n7840;
   wire n7835;
   wire n7831;
   wire n783;
   wire n7826;
   wire n7822;
   wire n7818;
   wire n7815;
   wire n7810;
   wire n7806;
   wire n7802;
   wire n7798;
   wire n7793;
   wire n779;
   wire n7788;
   wire n7784;
   wire n7779;
   wire n7776;
   wire n7773;
   wire n7768;
   wire n7764;
   wire n7760;
   wire n7756;
   wire n7751;
   wire n7746;
   wire n7741;
   wire n774;
   wire n7737;
   wire n7732;
   wire n7728;
   wire n7723;
   wire n7719;
   wire n7714;
   wire n7709;
   wire n7704;
   wire n7700;
   wire n770;
   wire n7695;
   wire n7691;
   wire n7686;
   wire n7681;
   wire n7676;
   wire n7671;
   wire n7666;
   wire n7661;
   wire n7658;
   wire n7654;
   wire n765;
   wire n7649;
   wire n7644;
   wire n7640;
   wire n7635;
   wire n7631;
   wire n7626;
   wire n7622;
   wire n7618;
   wire n7613;
   wire n761;
   wire n7608;
   wire n7604;
   wire n7599;
   wire n7596;
   wire n7591;
   wire n7586;
   wire n7581;
   wire n7577;
   wire n7572;
   wire n7567;
   wire n7563;
   wire n756;
   wire n7558;
   wire n7553;
   wire n7548;
   wire n7543;
   wire n7539;
   wire n7535;
   wire n7530;
   wire n7527;
   wire n7522;
   wire n7518;
   wire n7513;
   wire n751;
   wire n7509;
   wire n7505;
   wire n7501;
   wire n7496;
   wire n7492;
   wire n7487;
   wire n7482;
   wire n7478;
   wire n7473;
   wire n7468;
   wire n7463;
   wire n746;
   wire n7459;
   wire n7454;
   wire n7450;
   wire n7446;
   wire n7442;
   wire n7437;
   wire n7432;
   wire n7427;
   wire n7422;
   wire n7417;
   wire n7413;
   wire n741;
   wire n7408;
   wire n7404;
   wire n7400;
   wire n7395;
   wire n7391;
   wire n7386;
   wire n7381;
   wire n7376;
   wire n7372;
   wire n7368;
   wire n7363;
   wire n736;
   wire n7359;
   wire n7354;
   wire n7349;
   wire n7344;
   wire n7340;
   wire n7335;
   wire n7330;
   wire n7326;
   wire n7321;
   wire n732;
   wire n7316;
   wire n7312;
   wire n7307;
   wire n7302;
   wire n7297;
   wire n7292;
   wire n7288;
   wire n7284;
   wire n7280;
   wire n7275;
   wire n7270;
   wire n727;
   wire n7265;
   wire n7260;
   wire n7256;
   wire n7252;
   wire n7249;
   wire n7245;
   wire n7240;
   wire n7235;
   wire n7230;
   wire n7226;
   wire n7221;
   wire n722;
   wire n7216;
   wire n7212;
   wire n7207;
   wire n7203;
   wire n7199;
   wire n7194;
   wire n7190;
   wire n7185;
   wire n7182;
   wire n718;
   wire n7177;
   wire n7172;
   wire n7167;
   wire n7164;
   wire n7160;
   wire n7155;
   wire n7151;
   wire n7147;
   wire n7142;
   wire n7138;
   wire n7133;
   wire n713;
   wire n7128;
   wire n7125;
   wire n7120;
   wire n7116;
   wire n7111;
   wire n7107;
   wire n7102;
   wire n7098;
   wire n7093;
   wire n7089;
   wire n7085;
   wire n7082;
   wire n708;
   wire n7077;
   wire n7072;
   wire n7067;
   wire n7062;
   wire n7058;
   wire n7053;
   wire n7049;
   wire n7045;
   wire n7041;
   wire n7036;
   wire n7032;
   wire n703;
   wire n7027;
   wire n7023;
   wire n7018;
   wire n7013;
   wire n7009;
   wire n7005;
   wire n7000;
   wire n6995;
   wire n6990;
   wire n6986;
   wire n6982;
   wire n698;
   wire n6977;
   wire n6974;
   wire n6969;
   wire n6964;
   wire n6960;
   wire n6957;
   wire n6952;
   wire n6947;
   wire n6943;
   wire n6938;
   wire n6934;
   wire n693;
   wire n6929;
   wire n6924;
   wire n6919;
   wire n6915;
   wire n6910;
   wire n6906;
   wire n6902;
   wire n6899;
   wire n6895;
   wire n6890;
   wire n6886;
   wire n6881;
   wire n688;
   wire n6876;
   wire n6872;
   wire n6867;
   wire n6863;
   wire n6860;
   wire n6855;
   wire n6850;
   wire n6845;
   wire n6840;
   wire n6836;
   wire n6831;
   wire n683;
   wire n6826;
   wire n6822;
   wire n6818;
   wire n6813;
   wire n6809;
   wire n6806;
   wire n6801;
   wire n6796;
   wire n6793;
   wire n6788;
   wire n6783;
   wire n678;
   wire n6779;
   wire n6774;
   wire n6770;
   wire n6765;
   wire n6761;
   wire n6756;
   wire n6752;
   wire n6749;
   wire n6746;
   wire n6741;
   wire n6736;
   wire n6732;
   wire n673;
   wire n6727;
   wire n6722;
   wire n6717;
   wire n6713;
   wire n6709;
   wire n6704;
   wire n6700;
   wire n6695;
   wire n6691;
   wire n669;
   wire n6687;
   wire n6682;
   wire n6678;
   wire n6674;
   wire n6669;
   wire n6665;
   wire n6661;
   wire n6656;
   wire n6652;
   wire n6648;
   wire n6643;
   wire n664;
   wire n6638;
   wire n6634;
   wire n6629;
   wire n6624;
   wire n6619;
   wire n6615;
   wire n6611;
   wire n6606;
   wire n6601;
   wire n6596;
   wire n6591;
   wire n659;
   wire n6586;
   wire n6583;
   wire n6578;
   wire n6574;
   wire n6570;
   wire n6566;
   wire n6563;
   wire n6558;
   wire n6554;
   wire n6550;
   wire n6545;
   wire n6540;
   wire n654;
   wire n6535;
   wire n6531;
   wire n6527;
   wire n6522;
   wire n6519;
   wire n6515;
   wire n6511;
   wire n6507;
   wire n6502;
   wire n6498;
   wire n6493;
   wire n649;
   wire n6489;
   wire n6485;
   wire n6480;
   wire n6477;
   wire n6472;
   wire n6469;
   wire n6464;
   wire n6460;
   wire n6455;
   wire n6450;
   wire n6446;
   wire n6441;
   wire n644;
   wire n6437;
   wire n6432;
   wire n6427;
   wire n6423;
   wire n6419;
   wire n6415;
   wire n6411;
   wire n6407;
   wire n6403;
   wire n6399;
   wire n6395;
   wire n6390;
   wire n639;
   wire n6386;
   wire n6381;
   wire n6376;
   wire n6371;
   wire n6367;
   wire n6362;
   wire n6357;
   wire n6354;
   wire n6350;
   wire n6346;
   wire n6342;
   wire n634;
   wire n6337;
   wire n6332;
   wire n6329;
   wire n6324;
   wire n6319;
   wire n6316;
   wire n6311;
   wire n6306;
   wire n6302;
   wire n6299;
   wire n6294;
   wire n6290;
   wire n629;
   wire n6285;
   wire n6281;
   wire n6276;
   wire n6271;
   wire n6266;
   wire n6261;
   wire n6258;
   wire n6254;
   wire n625;
   wire n6249;
   wire n6244;
   wire n6239;
   wire n6235;
   wire n6231;
   wire n6227;
   wire n6222;
   wire n6218;
   wire n6214;
   wire n6209;
   wire n6204;
   wire n6200;
   wire n620;
   wire n6195;
   wire n6191;
   wire n6186;
   wire n6181;
   wire n6176;
   wire n6171;
   wire n6166;
   wire n6161;
   wire n6158;
   wire n6153;
   wire n615;
   wire n6148;
   wire n6145;
   wire n6140;
   wire n6136;
   wire n6132;
   wire n6128;
   wire n6124;
   wire n6119;
   wire n6114;
   wire n6110;
   wire n6106;
   wire n6102;
   wire n610;
   wire n6098;
   wire n6093;
   wire n6088;
   wire n6083;
   wire n6078;
   wire n6074;
   wire n6069;
   wire n6066;
   wire n6061;
   wire n6056;
   wire n6052;
   wire n605;
   wire n6047;
   wire n6043;
   wire n6038;
   wire n6034;
   wire n6029;
   wire n6024;
   wire n6019;
   wire n6014;
   wire n6009;
   wire n6006;
   wire n6002;
   wire n600;
   wire n5997;
   wire n5992;
   wire n5987;
   wire n5982;
   wire n5978;
   wire n5973;
   wire n5968;
   wire n5964;
   wire n5960;
   wire n5955;
   wire n5951;
   wire n595;
   wire n5947;
   wire n5943;
   wire n5938;
   wire n5934;
   wire n5930;
   wire n5925;
   wire n5920;
   wire n5917;
   wire n5912;
   wire n5908;
   wire n5903;
   wire n590;
   wire n5899;
   wire n5894;
   wire n5890;
   wire n5885;
   wire n5881;
   wire n5876;
   wire n5872;
   wire n5867;
   wire n5864;
   wire n5860;
   wire n5855;
   wire n5850;
   wire n585;
   wire n5845;
   wire n5840;
   wire n5836;
   wire n5833;
   wire n5828;
   wire n5824;
   wire n5819;
   wire n5814;
   wire n5809;
   wire n5805;
   wire n5801;
   wire n580;
   wire n5796;
   wire n5792;
   wire n5787;
   wire n5783;
   wire n5779;
   wire n5775;
   wire n5771;
   wire n5767;
   wire n5763;
   wire n576;
   wire n5758;
   wire n5753;
   wire n5748;
   wire n5744;
   wire n5739;
   wire n5735;
   wire n5731;
   wire n5727;
   wire n5722;
   wire n5717;
   wire n5713;
   wire n571;
   wire n5709;
   wire n5704;
   wire n5700;
   wire n5696;
   wire n5691;
   wire n5686;
   wire n5682;
   wire n5679;
   wire n5674;
   wire n5669;
   wire n5664;
   wire n5660;
   wire n566;
   wire n5655;
   wire n5651;
   wire n5648;
   wire n5643;
   wire n5638;
   wire n5633;
   wire n5628;
   wire n5623;
   wire n5618;
   wire n5613;
   wire n5610;
   wire n561;
   wire n5606;
   wire n5601;
   wire n5596;
   wire n5591;
   wire n5588;
   wire n5584;
   wire n5579;
   wire n5575;
   wire n5570;
   wire n5565;
   wire n5560;
   wire n556;
   wire n5556;
   wire n5552;
   wire n5547;
   wire n5543;
   wire n5539;
   wire n5534;
   wire n553;
   wire n5529;
   wire n5525;
   wire n5521;
   wire n5517;
   wire n5513;
   wire n5508;
   wire n5504;
   wire n5500;
   wire n5495;
   wire n5490;
   wire n5486;
   wire n5481;
   wire n548;
   wire n5477;
   wire n5472;
   wire n5469;
   wire n5464;
   wire n5460;
   wire n5455;
   wire n5451;
   wire n5446;
   wire n5441;
   wire n5437;
   wire n5433;
   wire n543;
   wire n5429;
   wire n5424;
   wire n5420;
   wire n5415;
   wire n5411;
   wire n5406;
   wire n5402;
   wire n5397;
   wire n5393;
   wire n5388;
   wire n5383;
   wire n5380;
   wire n538;
   wire n5375;
   wire n5370;
   wire n5366;
   wire n5362;
   wire n5358;
   wire n5353;
   wire n5349;
   wire n5344;
   wire n5339;
   wire n5335;
   wire n5330;
   wire n533;
   wire n5326;
   wire n5321;
   wire n5316;
   wire n5312;
   wire n5307;
   wire n5302;
   wire n5298;
   wire n5293;
   wire n5288;
   wire n5284;
   wire n528;
   wire n5279;
   wire n5274;
   wire n5269;
   wire n5265;
   wire n5261;
   wire n5256;
   wire n5251;
   wire n5246;
   wire n5242;
   wire n5239;
   wire n5234;
   wire n5230;
   wire n523;
   wire n5225;
   wire n5221;
   wire n5217;
   wire n5212;
   wire n5207;
   wire n5202;
   wire n5198;
   wire n5193;
   wire n5189;
   wire n5186;
   wire n5181;
   wire n518;
   wire n5178;
   wire n5173;
   wire n5169;
   wire n5164;
   wire n5159;
   wire n5156;
   wire n5151;
   wire n5148;
   wire n5143;
   wire n5139;
   wire n5134;
   wire n5130;
   wire n513;
   wire n5126;
   wire n5121;
   wire n5117;
   wire n5112;
   wire n5107;
   wire n5103;
   wire n5098;
   wire n5094;
   wire n5090;
   wire n5085;
   wire n5080;
   wire n508;
   wire n5075;
   wire n5070;
   wire n5066;
   wire n5061;
   wire n5056;
   wire n5053;
   wire n5048;
   wire n5045;
   wire n5040;
   wire n5035;
   wire n5031;
   wire n503;
   wire n5027;
   wire n5023;
   wire n5018;
   wire n5013;
   wire n5008;
   wire n5005;
   wire n5001;
   wire n4996;
   wire n4992;
   wire n4987;
   wire n4983;
   wire n498;
   wire n4979;
   wire n4974;
   wire n4969;
   wire n4965;
   wire n4961;
   wire n4957;
   wire n4952;
   wire n4947;
   wire n4944;
   wire n4940;
   wire n4936;
   wire n4931;
   wire n493;
   wire n4927;
   wire n4922;
   wire n4917;
   wire n4913;
   wire n4908;
   wire n4904;
   wire n4899;
   wire n4895;
   wire n4890;
   wire n4886;
   wire n4881;
   wire n488;
   wire n4877;
   wire n4872;
   wire n4867;
   wire n4862;
   wire n4857;
   wire n4853;
   wire n4848;
   wire n4843;
   wire n484;
   wire n4838;
   wire n4834;
   wire n4831;
   wire n4827;
   wire n4822;
   wire n4818;
   wire n4814;
   wire n4809;
   wire n4805;
   wire n4800;
   wire n4795;
   wire n4791;
   wire n479;
   wire n4787;
   wire n4782;
   wire n4778;
   wire n4774;
   wire n4769;
   wire n4765;
   wire n4760;
   wire n4755;
   wire n4750;
   wire n4745;
   wire n4742;
   wire n474;
   wire n4737;
   wire n4732;
   wire n4727;
   wire n4722;
   wire n4717;
   wire n4713;
   wire n4708;
   wire n4703;
   wire n470;
   wire n4699;
   wire n4694;
   wire n4690;
   wire n4686;
   wire n4681;
   wire n4678;
   wire n4673;
   wire n4669;
   wire n4665;
   wire n4660;
   wire n4656;
   wire n4651;
   wire n465;
   wire n4646;
   wire n4641;
   wire n4636;
   wire n4631;
   wire n4627;
   wire n4622;
   wire n4617;
   wire n4613;
   wire n4609;
   wire n4604;
   wire n4600;
   wire n460;
   wire n4596;
   wire n4591;
   wire n4586;
   wire n4581;
   wire n4577;
   wire n4572;
   wire n4567;
   wire n4562;
   wire n4558;
   wire n4553;
   wire n455;
   wire n4548;
   wire n4544;
   wire n4539;
   wire n4534;
   wire n4529;
   wire n4524;
   wire n4520;
   wire n4515;
   wire n4510;
   wire n451;
   wire n4505;
   wire n4501;
   wire n4496;
   wire n4491;
   wire n4487;
   wire n4482;
   wire n4478;
   wire n4473;
   wire n447;
   wire n4469;
   wire n4464;
   wire n4459;
   wire n4456;
   wire n4451;
   wire n4448;
   wire n4443;
   wire n4438;
   wire n4433;
   wire n443;
   wire n4428;
   wire n4424;
   wire n4419;
   wire n4414;
   wire n4410;
   wire n4405;
   wire n4401;
   wire n4397;
   wire n4392;
   wire n4388;
   wire n4384;
   wire n438;
   wire n4379;
   wire n4374;
   wire n4370;
   wire n4365;
   wire n4362;
   wire n4357;
   wire n4352;
   wire n4348;
   wire n4343;
   wire n434;
   wire n4338;
   wire n4333;
   wire n4330;
   wire n4326;
   wire n4322;
   wire n4318;
   wire n4313;
   wire n4309;
   wire n4304;
   wire n4299;
   wire n4294;
   wire n429;
   wire n4289;
   wire n4284;
   wire n4280;
   wire n4276;
   wire n4271;
   wire n4267;
   wire n4263;
   wire n4258;
   wire n4253;
   wire n4249;
   wire n4245;
   wire n4240;
   wire n424;
   wire n4235;
   wire n4231;
   wire n4226;
   wire n4221;
   wire n4217;
   wire n4212;
   wire n4207;
   wire n4203;
   wire n420;
   wire n4199;
   wire n4194;
   wire n4191;
   wire n4186;
   wire n4181;
   wire n4176;
   wire n4171;
   wire n4166;
   wire n4161;
   wire n4158;
   wire n4153;
   wire n415;
   wire n4148;
   wire n4145;
   wire n4140;
   wire n4135;
   wire n4131;
   wire n4126;
   wire n4121;
   wire n4116;
   wire n4112;
   wire n4107;
   wire n4102;
   wire n410;
   wire n4098;
   wire n4094;
   wire n4089;
   wire n4084;
   wire n4079;
   wire n4075;
   wire n4071;
   wire n4068;
   wire n4063;
   wire n4059;
   wire n4055;
   wire n4051;
   wire n405;
   wire n4046;
   wire n4042;
   wire n4037;
   wire n4033;
   wire n4029;
   wire n4024;
   wire n4020;
   wire n4016;
   wire n4011;
   wire n4007;
   wire n4002;
   wire n400;
   wire n3998;
   wire n3993;
   wire n3989;
   wire n3985;
   wire n3981;
   wire n3976;
   wire n3972;
   wire n3967;
   wire n3962;
   wire n3957;
   wire n3953;
   wire n395;
   wire n3949;
   wire n3945;
   wire n3941;
   wire n3936;
   wire n3932;
   wire n3927;
   wire n3922;
   wire n3917;
   wire n3913;
   wire n3908;
   wire n3904;
   wire n390;
   wire n3899;
   wire n3896;
   wire n3891;
   wire n3886;
   wire n3881;
   wire n3877;
   wire n3872;
   wire n3867;
   wire n3864;
   wire n3859;
   wire n3855;
   wire n3851;
   wire n385;
   wire n3846;
   wire n3841;
   wire n3836;
   wire n3831;
   wire n3827;
   wire n3822;
   wire n3817;
   wire n3813;
   wire n3809;
   wire n3805;
   wire n3801;
   wire n380;
   wire n3796;
   wire n3791;
   wire n3787;
   wire n3782;
   wire n3777;
   wire n3773;
   wire n3770;
   wire n3765;
   wire n3761;
   wire n3756;
   wire n3752;
   wire n375;
   wire n3747;
   wire n3742;
   wire n3737;
   wire n3733;
   wire n3729;
   wire n3725;
   wire n3720;
   wire n3716;
   wire n3711;
   wire n3707;
   wire n3703;
   wire n370;
   wire n3698;
   wire n3693;
   wire n3689;
   wire n3684;
   wire n3679;
   wire n3675;
   wire n3670;
   wire n3666;
   wire n3661;
   wire n366;
   wire n3658;
   wire n3655;
   wire n3651;
   wire n3647;
   wire n3642;
   wire n3638;
   wire n3633;
   wire n3628;
   wire n3623;
   wire n3618;
   wire n3614;
   wire n361;
   wire n3609;
   wire n3604;
   wire n3600;
   wire n3595;
   wire n3590;
   wire n3587;
   wire n3582;
   wire n3577;
   wire n3572;
   wire n357;
   wire n3567;
   wire n3564;
   wire n3559;
   wire n3555;
   wire n3551;
   wire n3546;
   wire n3542;
   wire n3537;
   wire n3532;
   wire n3528;
   wire n3524;
   wire n3520;
   wire n352;
   wire n3516;
   wire n3511;
   wire n3507;
   wire n3502;
   wire n3497;
   wire n3494;
   wire n349;
   wire n3489;
   wire n3484;
   wire n3479;
   wire n3474;
   wire n3469;
   wire n3464;
   wire n3459;
   wire n3455;
   wire n3450;
   wire n3445;
   wire n3440;
   wire n344;
   wire n3436;
   wire n3431;
   wire n3427;
   wire n3422;
   wire n3418;
   wire n3413;
   wire n3408;
   wire n3404;
   wire n3400;
   wire n3395;
   wire n3390;
   wire n339;
   wire n3386;
   wire n3383;
   wire n3379;
   wire n3374;
   wire n3370;
   wire n3365;
   wire n3361;
   wire n3356;
   wire n3352;
   wire n3348;
   wire n3343;
   wire n334;
   wire n3338;
   wire n3333;
   wire n3330;
   wire n3325;
   wire n3322;
   wire n3318;
   wire n3313;
   wire n3308;
   wire n3303;
   wire n3299;
   wire n3294;
   wire n3290;
   wire n329;
   wire n3285;
   wire n3280;
   wire n3276;
   wire n3272;
   wire n3268;
   wire n3263;
   wire n3258;
   wire n3254;
   wire n3249;
   wire n3244;
   wire n3240;
   wire n324;
   wire n3235;
   wire n3231;
   wire n3226;
   wire n3222;
   wire n3217;
   wire n3212;
   wire n3207;
   wire n3203;
   wire n3199;
   wire n3194;
   wire n3190;
   wire n319;
   wire n3186;
   wire n3182;
   wire n3178;
   wire n3174;
   wire n3170;
   wire n3165;
   wire n3162;
   wire n3157;
   wire n3152;
   wire n3148;
   wire n3143;
   wire n314;
   wire n3139;
   wire n3134;
   wire n3130;
   wire n3126;
   wire n3121;
   wire n3117;
   wire n3114;
   wire n3110;
   wire n3105;
   wire n3102;
   wire n310;
   wire n3097;
   wire n3092;
   wire n3087;
   wire n3082;
   wire n3078;
   wire n3074;
   wire n3069;
   wire n3065;
   wire n3061;
   wire n3056;
   wire n3052;
   wire n305;
   wire n3047;
   wire n3042;
   wire n3037;
   wire n3033;
   wire n3030;
   wire n3025;
   wire n3020;
   wire n3015;
   wire n3010;
   wire n3005;
   wire n3000;
   wire n300;
   wire n2996;
   wire n2991;
   wire n2986;
   wire n2981;
   wire n2976;
   wire n2972;
   wire n2967;
   wire n2963;
   wire n2958;
   wire n2953;
   wire n295;
   wire n2948;
   wire n2944;
   wire n2939;
   wire n2935;
   wire n2930;
   wire n2926;
   wire n2922;
   wire n2918;
   wire n2913;
   wire n291;
   wire n2908;
   wire n2904;
   wire n2900;
   wire n2895;
   wire n2890;
   wire n2885;
   wire n2882;
   wire n2877;
   wire n2873;
   wire n2869;
   wire n2864;
   wire n2860;
   wire n286;
   wire n2855;
   wire n2850;
   wire n2845;
   wire n2840;
   wire n2836;
   wire n2831;
   wire n2827;
   wire n2823;
   wire n2819;
   wire n2814;
   wire n2810;
   wire n281;
   wire n2805;
   wire n2801;
   wire n2797;
   wire n2792;
   wire n2788;
   wire n2784;
   wire n2781;
   wire n2776;
   wire n2771;
   wire n2767;
   wire n2762;
   wire n276;
   wire n2758;
   wire n2753;
   wire n2748;
   wire n2745;
   wire n2741;
   wire n2737;
   wire n2732;
   wire n2727;
   wire n2723;
   wire n2718;
   wire n2713;
   wire n271;
   wire n2709;
   wire n2705;
   wire n2701;
   wire n2696;
   wire n2692;
   wire n2687;
   wire n2682;
   wire n2679;
   wire n2675;
   wire n2670;
   wire n2665;
   wire n2660;
   wire n266;
   wire n2656;
   wire n2651;
   wire n2647;
   wire n2642;
   wire n2637;
   wire n2632;
   wire n2627;
   wire n2622;
   wire n2618;
   wire n2615;
   wire n2610;
   wire n2605;
   wire n2601;
   wire n2597;
   wire n2594;
   wire n2590;
   wire n2585;
   wire n2580;
   wire n2575;
   wire n2570;
   wire n2566;
   wire n2561;
   wire n2556;
   wire n2552;
   wire n2547;
   wire n2543;
   wire n2539;
   wire n2534;
   wire n2529;
   wire n2524;
   wire n2519;
   wire n2515;
   wire n2510;
   wire n2505;
   wire n2500;
   wire n2496;
   wire n2493;
   wire n2488;
   wire n2484;
   wire n2479;
   wire n2474;
   wire n2470;
   wire n2465;
   wire n2462;
   wire n2457;
   wire n2452;
   wire n2448;
   wire n2444;
   wire n2440;
   wire n2435;
   wire n2430;
   wire n2426;
   wire n2422;
   wire n2417;
   wire n2414;
   wire n2409;
   wire n2404;
   wire n2399;
   wire n2395;
   wire n2391;
   wire n2386;
   wire n2381;
   wire n2377;
   wire n2373;
   wire n2370;
   wire n2365;
   wire n2360;
   wire n2355;
   wire n2350;
   wire n2347;
   wire n2342;
   wire n2338;
   wire n2334;
   wire n2329;
   wire n2324;
   wire n2321;
   wire n2316;
   wire n2312;
   wire n2307;
   wire n2303;
   wire n2298;
   wire n2293;
   wire n2288;
   wire n2284;
   wire n2280;
   wire n2275;
   wire n2270;
   wire n2265;
   wire n2260;
   wire n2256;
   wire n2251;
   wire n2247;
   wire n2242;
   wire n2237;
   wire n2232;
   wire n2227;
   wire n2222;
   wire n2218;
   wire n2213;
   wire n2208;
   wire n2203;
   wire n2199;
   wire n2194;
   wire n2189;
   wire n2186;
   wire n2181;
   wire n2177;
   wire n2172;
   wire n2167;
   wire n2162;
   wire n2157;
   wire n2152;
   wire n2149;
   wire n2144;
   wire n2140;
   wire n2136;
   wire n2132;
   wire n2127;
   wire n2122;
   wire n2119;
   wire n2115;
   wire n2111;
   wire n2106;
   wire n2102;
   wire n2098;
   wire n2093;
   wire n2088;
   wire n2084;
   wire n2079;
   wire n2074;
   wire n2070;
   wire n2065;
   wire n2060;
   wire n2055;
   wire n2051;
   wire n2046;
   wire n2041;
   wire n2036;
   wire n2031;
   wire n2026;
   wire n2021;
   wire n2016;
   wire n2011;
   wire n2007;
   wire n2002;
   wire n1998;
   wire n1993;
   wire n1988;
   wire n1983;
   wire n1978;
   wire n1973;
   wire n1969;
   wire n1964;
   wire n1959;
   wire n1954;
   wire n1950;
   wire n1945;
   wire n1941;
   wire n1936;
   wire n1932;
   wire n1927;
   wire n1922;
   wire n1918;
   wire n1913;
   wire n1908;
   wire n1903;
   wire n1898;
   wire n1893;
   wire n1888;
   wire n1883;
   wire n1878;
   wire n1874;
   wire n1869;
   wire n1865;
   wire n1860;
   wire n1855;
   wire n1851;
   wire n1846;
   wire n1841;
   wire n1836;
   wire n1832;
   wire n1827;
   wire n1822;
   wire n1817;
   wire n1812;
   wire n1807;
   wire n1802;
   wire n1797;
   wire n1792;
   wire n1787;
   wire n1782;
   wire n1779;
   wire n1775;
   wire n1770;
   wire n1765;
   wire n1761;
   wire n1756;
   wire n1752;
   wire n1747;
   wire n1742;
   wire n1737;
   wire n1732;
   wire n1727;
   wire n1722;
   wire n1718;
   wire n1714;
   wire n1709;
   wire n1704;
   wire n1701;
   wire n1696;
   wire n1691;
   wire n1686;
   wire n1681;
   wire n1677;
   wire n1673;
   wire n1668;
   wire n1663;
   wire n1658;
   wire n1653;
   wire n1649;
   wire n1644;
   wire n1639;
   wire n1634;
   wire n1629;
   wire n1624;
   wire n1619;
   wire n1615;
   wire n1610;
   wire n1605;
   wire n1600;
   wire n1596;
   wire n1591;
   wire n1587;
   wire n1582;
   wire n1577;
   wire n1572;
   wire n1568;
   wire n1564;
   wire n1560;
   wire n1555;
   wire n1551;
   wire n1546;
   wire n1542;
   wire n1538;
   wire n1533;
   wire n1528;
   wire n1524;
   wire n1519;
   wire n1515;
   wire n1510;
   wire n1506;
   wire n1501;
   wire n1496;
   wire n1491;
   wire n1487;
   wire n1482;
   wire n1478;
   wire n1474;
   wire n1469;
   wire n1465;
   wire n1460;
   wire n1455;
   wire n1451;
   wire n1446;
   wire n1442;
   wire n1438;
   wire n1433;
   wire n1428;
   wire n1423;
   wire n1419;
   wire n1414;
   wire n1410;
   wire n1405;
   wire n1400;
   wire n1396;
   wire n1391;
   wire n1386;
   wire n1383;
   wire n1378;
   wire n1373;
   wire n1368;
   wire n1363;
   wire n1359;
   wire n1355;
   wire n1350;
   wire n1345;
   wire n1340;
   wire n1335;
   wire n1331;
   wire n1326;
   wire n1322;
   wire n1318;
   wire n1314;
   wire n1309;
   wire n1305;
   wire n1300;
   wire n1295;
   wire n1291;
   wire n1287;
   wire n1282;
   wire n1277;
   wire n1272;
   wire n1267;
   wire n1262;
   wire n1258;
   wire n1253;
   wire n1248;
   wire n1244;
   wire n1240;
   wire n1236;
   wire n1232;
   wire n1228;
   wire n1224;
   wire n1219;
   wire n1214;
   wire n1210;
   wire n1205;
   wire n1200;
   wire n1195;
   wire n1191;
   wire n1187;
   wire n1183;
   wire n1178;
   wire n1173;
   wire n1168;
   wire n1163;
   wire n1158;
   wire n1153;
   wire n1148;
   wire n1144;
   wire n1140;
   wire n1135;
   wire n1130;
   wire n1125;
   wire n1121;
   wire n1116;
   wire n1111;
   wire n1106;
   wire n1102;
   wire n1097;
   wire n1093;
   wire n1089;
   wire n1085;
   wire n1081;
   wire n1077;
   wire n1072;
   wire n1067;
   wire n1062;
   wire n1058;
   wire n1053;
   wire n1049;
   wire n1044;
   wire n1039;
   wire n1034;
   wire n1029;
   wire n1024;
   wire n1020;
   wire n10158;
   wire n10154;
   wire n10150;
   wire n1015;
   wire n10145;
   wire n10141;
   wire n10137;
   wire n10132;
   wire n10128;
   wire n10124;
   wire n10120;
   wire n10116;
   wire n10112;
   wire n10107;
   wire n10103;
   wire n1010;
   wire n10099;
   wire n10094;
   wire n10089;
   wire n10084;
   wire n10079;
   wire n10074;
   wire n10070;
   wire n10066;
   wire n10061;
   wire n10056;
   wire n10052;
   wire n1005;
   wire n10047;
   wire n10042;
   wire n10037;
   wire n10032;
   wire n10028;
   wire n10023;
   wire n10019;
   wire n10014;
   wire n10010;
   wire n10006;
   wire n10001;
   wire n1000;
   wire clk;
   wire _net_7824;
   wire _net_7823;
   wire _net_7822;
   wire _net_7821;
   wire _net_7820;
   wire _net_7819;
   wire _net_7818;
   wire _net_7817;
   wire _net_7816;
   wire _net_7815;
   wire _net_7814;
   wire _net_7813;
   wire _net_7812;
   wire _net_7811;
   wire _net_7810;
   wire _net_7809;
   wire _net_7808;
   wire _net_7806;
   wire _net_7805;
   wire _net_7804;
   wire _net_7803;
   wire _net_7801;
   wire _net_7800;
   wire _net_7798;
   wire _net_7797;
   wire _net_7796;
   wire _net_7795;
   wire _net_7794;
   wire _net_7793;
   wire _net_7791;
   wire _net_7789;
   wire _net_7788;
   wire _net_7787;
   wire _net_7786;
   wire _net_7785;
   wire _net_7784;
   wire _net_7783;
   wire _net_7782;
   wire _net_7781;
   wire _net_7768;
   wire _net_7765;
   wire _net_7763;
   wire _net_7761;
   wire _net_7759;
   wire _net_7757;
   wire _net_7755;
   wire _net_7753;
   wire _net_7751;
   wire _net_7749;
   wire _net_7748;
   wire _net_7747;
   wire _net_7746;
   wire _net_7745;
   wire _net_7736;
   wire _net_7735;
   wire _net_7734;
   wire _net_7733;
   wire _net_7732;
   wire _net_7731;
   wire _net_7730;
   wire _net_7729;
   wire _net_7728;
   wire _net_7727;
   wire _net_7726;
   wire _net_7725;
   wire _net_7724;
   wire _net_7723;
   wire _net_7722;
   wire _net_7721;
   wire _net_7720;
   wire _net_7719;
   wire _net_7718;
   wire _net_7717;
   wire _net_7716;
   wire _net_7707;
   wire _net_7706;
   wire _net_7705;
   wire _net_7704;
   wire _net_7703;
   wire _net_7702;
   wire _net_7701;
   wire _net_7700;
   wire _net_7699;
   wire _net_7698;
   wire _net_7697;
   wire _net_7696;
   wire _net_7695;
   wire _net_7694;
   wire _net_7693;
   wire _net_7692;
   wire _net_7690;
   wire _net_7689;
   wire _net_7688;
   wire _net_7687;
   wire _net_7686;
   wire _net_7685;
   wire _net_7684;
   wire _net_7683;
   wire _net_7682;
   wire _net_7681;
   wire _net_7667;
   wire _net_7666;
   wire _net_7665;
   wire _net_7664;
   wire _net_7663;
   wire _net_7662;
   wire _net_7661;
   wire _net_7660;
   wire _net_7659;
   wire _net_7658;
   wire _net_7657;
   wire _net_7656;
   wire _net_7655;
   wire _net_7654;
   wire _net_7653;
   wire _net_7652;
   wire _net_7651;
   wire _net_7650;
   wire _net_7649;
   wire _net_7648;
   wire _net_7635;
   wire _net_7634;
   wire _net_7633;
   wire _net_7632;
   wire _net_7631;
   wire _net_7630;
   wire _net_7629;
   wire _net_7628;
   wire _net_7627;
   wire _net_7626;
   wire _net_7625;
   wire _net_7624;
   wire _net_7623;
   wire _net_7622;
   wire _net_7621;
   wire _net_7620;
   wire _net_7619;
   wire _net_7618;
   wire _net_7617;
   wire _net_7616;
   wire _net_7603;
   wire _net_7602;
   wire _net_7601;
   wire _net_7600;
   wire _net_7599;
   wire _net_7598;
   wire _net_7597;
   wire _net_7596;
   wire _net_7595;
   wire _net_7594;
   wire _net_7593;
   wire _net_7592;
   wire _net_7591;
   wire _net_7590;
   wire _net_7589;
   wire _net_7588;
   wire _net_7587;
   wire _net_7586;
   wire _net_7585;
   wire _net_7584;
   wire _net_7583;
   wire _net_7582;
   wire _net_7581;
   wire _net_7580;
   wire _net_7579;
   wire _net_7578;
   wire _net_7577;
   wire _net_7576;
   wire _net_7575;
   wire _net_7574;
   wire _net_7573;
   wire _net_7572;
   wire _net_7571;
   wire _net_7570;
   wire _net_7569;
   wire _net_7568;
   wire _net_7567;
   wire _net_7566;
   wire _net_7565;
   wire _net_7564;
   wire _net_7563;
   wire _net_7562;
   wire _net_7561;
   wire _net_7560;
   wire _net_7559;
   wire _net_7558;
   wire _net_7557;
   wire _net_7556;
   wire _net_7555;
   wire _net_7554;
   wire _net_7553;
   wire _net_7552;
   wire _net_7535;
   wire _net_7534;
   wire _net_7533;
   wire _net_7532;
   wire _net_7531;
   wire _net_7530;
   wire _net_7516;
   wire _net_7515;
   wire _net_7514;
   wire _net_7513;
   wire _net_7512;
   wire _net_7511;
   wire _net_7510;
   wire _net_7509;
   wire _net_7508;
   wire _net_7507;
   wire _net_7506;
   wire _net_7505;
   wire _net_7504;
   wire _net_7503;
   wire _net_7502;
   wire _net_7501;
   wire _net_7500;
   wire _net_7499;
   wire _net_7498;
   wire _net_7497;
   wire _net_7484;
   wire _net_7483;
   wire _net_7482;
   wire _net_7481;
   wire _net_7480;
   wire _net_7479;
   wire _net_7478;
   wire _net_7477;
   wire _net_7476;
   wire _net_7475;
   wire _net_7474;
   wire _net_7473;
   wire _net_7472;
   wire _net_7471;
   wire _net_7470;
   wire _net_7469;
   wire _net_7468;
   wire _net_7467;
   wire _net_7466;
   wire _net_7465;
   wire _net_7452;
   wire _net_7451;
   wire _net_7450;
   wire _net_7449;
   wire _net_7448;
   wire _net_7447;
   wire _net_7446;
   wire _net_7445;
   wire _net_7444;
   wire _net_7443;
   wire _net_7442;
   wire _net_7441;
   wire _net_7440;
   wire _net_7439;
   wire _net_7438;
   wire _net_7437;
   wire _net_7436;
   wire _net_7435;
   wire _net_7434;
   wire _net_7433;
   wire _net_7432;
   wire _net_7431;
   wire _net_7430;
   wire _net_7429;
   wire _net_7428;
   wire _net_7427;
   wire _net_7426;
   wire _net_7425;
   wire _net_7424;
   wire _net_7423;
   wire _net_7422;
   wire _net_7421;
   wire _net_7420;
   wire _net_7419;
   wire _net_7418;
   wire _net_7417;
   wire _net_7416;
   wire _net_7415;
   wire _net_7414;
   wire _net_7413;
   wire _net_7412;
   wire _net_7411;
   wire _net_7410;
   wire _net_7409;
   wire _net_7408;
   wire _net_7407;
   wire _net_7406;
   wire _net_7405;
   wire _net_7404;
   wire _net_7403;
   wire _net_7402;
   wire _net_7401;
   wire _net_7384;
   wire _net_7383;
   wire _net_7382;
   wire _net_7381;
   wire _net_7380;
   wire _net_7379;
   wire _net_7365;
   wire _net_7364;
   wire _net_7363;
   wire _net_7362;
   wire _net_7361;
   wire _net_7360;
   wire _net_7359;
   wire _net_7358;
   wire _net_7357;
   wire _net_7356;
   wire _net_7355;
   wire _net_7354;
   wire _net_7353;
   wire _net_7352;
   wire _net_7351;
   wire _net_7350;
   wire _net_7349;
   wire _net_7348;
   wire _net_7347;
   wire _net_7346;
   wire _net_7333;
   wire _net_7332;
   wire _net_7331;
   wire _net_7330;
   wire _net_7329;
   wire _net_7328;
   wire _net_7327;
   wire _net_7326;
   wire _net_7325;
   wire _net_7324;
   wire _net_7323;
   wire _net_7322;
   wire _net_7321;
   wire _net_7320;
   wire _net_7319;
   wire _net_7318;
   wire _net_7317;
   wire _net_7316;
   wire _net_7315;
   wire _net_7314;
   wire _net_7301;
   wire _net_7300;
   wire _net_7299;
   wire _net_7298;
   wire _net_7297;
   wire _net_7296;
   wire _net_7295;
   wire _net_7294;
   wire _net_7293;
   wire _net_7292;
   wire _net_7291;
   wire _net_7290;
   wire _net_7289;
   wire _net_7288;
   wire _net_7287;
   wire _net_7286;
   wire _net_7285;
   wire _net_7284;
   wire _net_7283;
   wire _net_7282;
   wire _net_7281;
   wire _net_7280;
   wire _net_7279;
   wire _net_7278;
   wire _net_7277;
   wire _net_7276;
   wire _net_7275;
   wire _net_7274;
   wire _net_7273;
   wire _net_7272;
   wire _net_7271;
   wire _net_7270;
   wire _net_7269;
   wire _net_7268;
   wire _net_7267;
   wire _net_7266;
   wire _net_7265;
   wire _net_7264;
   wire _net_7263;
   wire _net_7262;
   wire _net_7261;
   wire _net_7260;
   wire _net_7259;
   wire _net_7258;
   wire _net_7257;
   wire _net_7256;
   wire _net_7255;
   wire _net_7254;
   wire _net_7253;
   wire _net_7252;
   wire _net_7251;
   wire _net_7250;
   wire _net_7233;
   wire _net_7232;
   wire _net_7230;
   wire _net_7229;
   wire _net_7228;
   wire _net_7227;
   wire _net_7098;
   wire _net_7097;
   wire _net_7095;
   wire _net_7094;
   wire _net_7093;
   wire _net_7092;
   wire _net_6963;
   wire _net_6962;
   wire _net_6960;
   wire _net_6959;
   wire _net_6958;
   wire _net_6957;
   wire _net_6828;
   wire _net_6827;
   wire _net_6825;
   wire _net_6824;
   wire _net_6823;
   wire _net_6822;
   wire _net_6693;
   wire _net_6692;
   wire _net_6690;
   wire _net_6689;
   wire _net_6688;
   wire _net_6687;
   wire _net_6558;
   wire _net_6557;
   wire _net_6555;
   wire _net_6554;
   wire _net_6553;
   wire _net_6552;
   wire _net_6423;
   wire _net_6422;
   wire _net_6421;
   wire _net_6420;
   wire _net_6419;
   wire _net_6418;
   wire _net_6415;
   wire _net_6414;
   wire _net_6413;
   wire _net_6411;
   wire _net_6410;
   wire _net_6409;
   wire _net_6408;
   wire _net_6407;
   wire _net_6406;
   wire _net_6405;
   wire _net_6404;
   wire _net_6402;
   wire _net_6401;
   wire _net_6319;
   wire _net_6298;
   wire _net_6297;
   wire _net_6296;
   wire _net_6295;
   wire _net_6294;
   wire _net_6293;
   wire _net_6292;
   wire _net_6291;
   wire _net_6290;
   wire _net_6289;
   wire _net_6288;
   wire _net_6287;
   wire _net_6286;
   wire _net_6285;
   wire _net_6284;
   wire _net_6283;
   wire _net_6282;
   wire _net_6281;
   wire _net_6280;
   wire _net_6259;
   wire _net_6239;
   wire _net_6222;
   wire _net_6221;
   wire _net_6220;
   wire _net_6219;
   wire _net_6210;
   wire _net_6209;
   wire _net_6208;
   wire _net_6207;
   wire _net_6206;
   wire _net_6205;
   wire _net_6204;
   wire _net_6203;
   wire _net_6202;
   wire _net_6201;
   wire _net_6200;
   wire _net_6199;
   wire _net_6194;
   wire _net_6189;
   wire _net_6188;
   wire _net_6187;
   wire _net_6186;
   wire _net_6185;
   wire _net_6184;
   wire _net_6183;
   wire _net_6182;
   wire _net_6181;
   wire _net_6180;
   wire _net_6179;
   wire _net_6178;
   wire _net_6177;
   wire _net_6176;
   wire _net_6175;
   wire _net_6174;
   wire _net_6173;
   wire _net_6172;
   wire _net_6171;
   wire _net_6170;
   wire _net_6169;
   wire _net_6168;
   wire _net_6167;
   wire _net_6166;
   wire _net_6165;
   wire _net_6164;
   wire _net_6163;
   wire _net_6162;
   wire _net_6161;
   wire _net_6160;
   wire _net_6159;
   wire _net_6158;
   wire _net_6157;
   wire _net_6156;
   wire _net_6155;
   wire _net_6154;
   wire _net_6153;
   wire _net_6152;
   wire _net_6151;
   wire _net_6150;
   wire _net_6149;
   wire _net_6148;
   wire _net_6147;
   wire _net_6146;
   wire _net_6145;
   wire _net_6144;
   wire _net_6143;
   wire _net_6142;
   wire _net_6141;
   wire _net_6140;
   wire _net_6139;
   wire _net_6138;
   wire _net_6137;
   wire _net_6136;
   wire _net_6135;
   wire _net_6134;
   wire _net_6133;
   wire _net_6132;
   wire _net_6131;
   wire _net_6130;
   wire _net_6129;
   wire _net_6128;
   wire _net_6127;
   wire _net_6126;
   wire _net_6125;
   wire _net_6124;
   wire _net_6123;
   wire _net_6122;
   wire _net_6121;
   wire _net_6120;
   wire _net_6119;
   wire _net_6118;
   wire _net_6117;
   wire _net_6116;
   wire _net_6115;
   wire _net_6114;
   wire _net_6113;
   wire _net_6112;
   wire _net_6111;
   wire _net_6110;
   wire _net_6109;
   wire _net_6108;
   wire _net_6107;
   wire _net_6106;
   wire _net_6105;
   wire _net_6104;
   wire _net_6103;
   wire _net_6102;
   wire _net_6101;
   wire _net_6100;
   wire _net_6099;
   wire _net_6098;
   wire _net_6097;
   wire _net_6096;
   wire _net_6095;
   wire _net_6094;
   wire _net_6093;
   wire _net_6092;
   wire _net_6091;
   wire _net_6090;
   wire _net_6089;
   wire _net_6088;
   wire _net_6087;
   wire _net_6086;
   wire _net_6085;
   wire _net_6084;
   wire _net_6083;
   wire _net_6082;
   wire _net_6081;
   wire _net_6080;
   wire _net_6079;
   wire _net_6078;
   wire _net_6077;
   wire _net_6076;
   wire _net_6075;
   wire _net_6074;
   wire _net_6073;
   wire _net_6072;
   wire _net_6071;
   wire _net_6070;
   wire _net_6069;
   wire _net_6068;
   wire _net_6067;
   wire _net_6066;
   wire _net_6065;
   wire _net_6064;
   wire _net_6063;
   wire _net_6062;
   wire _net_6052;
   wire _net_6051;
   wire _net_6050;
   wire _net_6049;
   wire _net_6048;
   wire _net_6045;
   wire _net_6044;
   wire _net_6043;
   wire _net_6042;
   wire _net_6041;
   wire _net_6040;
   wire _net_6039;
   wire _net_6038;
   wire _net_6037;
   wire _net_6034;
   wire _net_6033;
   wire _net_6032;
   wire _net_6031;
   wire _net_6030;
   wire _net_6029;
   wire _net_6028;
   wire _net_6027;
   wire _net_6026;
   wire _net_6023;
   wire _net_6022;
   wire _net_6021;
   wire _net_6020;
   wire _net_6019;
   wire _net_6018;
   wire _net_6017;
   wire _net_6016;
   wire _net_6015;
   wire _net_6012;
   wire _net_6011;
   wire _net_6010;
   wire _net_6009;
   wire _net_6008;
   wire _net_6007;
   wire _net_6006;
   wire _net_6005;
   wire _net_6004;
   wire _net_6002;
   wire _net_6001;
   wire _net_6000;
   wire _net_5999;
   wire _net_5998;
   wire _net_5997;
   wire _net_5996;
   wire _net_5995;
   wire _net_5994;
   wire _net_5993;
   wire _net_5991;
   wire _net_5990;
   wire _net_5989;
   wire _net_5988;
   wire _net_5987;
   wire _net_5986;
   wire _net_5985;
   wire _net_5984;
   wire _net_5983;
   wire _net_5982;
   wire _net_5981;
   wire _net_5980;
   wire _net_5979;
   wire _net_5978;
   wire _net_5977;
   wire _net_5976;
   wire _net_5975;
   wire _net_5974;
   wire _net_5973;
   wire _net_5972;
   wire _net_5971;
   wire _net_5970;
   wire _net_5969;
   wire _net_5968;
   wire _net_5967;
   wire _net_5966;
   wire _net_5965;
   wire _net_5964;
   wire _net_5963;
   wire _net_5962;
   wire _net_5961;
   wire _net_5960;
   wire _net_5924;
   wire _net_5922;
   wire _net_5920;
   wire _net_5859;
   wire _net_5857;
   wire _net_5856;
   wire _net_5855;
   wire _net_5854;
   wire _net_5853;
   wire _net_5852;
   wire _net_5851;
   wire _net_5850;
   wire _net_5848;
   wire _net_392;
   wire _net_299;
   wire _net_298;
   wire _net_295;
   wire _net_294;
   wire _net_293;
   wire _net_292;
   wire _net_291;
   wire _net_290;
   wire _net_289;
   wire _net_288;
   wire _net_287;
   wire _net_284;
   wire _net_283;
   wire _net_282;
   wire _net_281;
   wire _net_280;
   wire _net_279;
   wire _net_278;
   wire _net_277;
   wire _net_276;
   wire _net_273;
   wire _net_272;
   wire _net_271;
   wire _net_270;
   wire _net_269;
   wire _net_268;
   wire _net_267;
   wire _net_266;
   wire _net_265;
   wire _net_264;
   wire _net_263;
   wire _net_262;
   wire _net_229;
   wire _net_228;
   wire _net_227;
   wire _net_226;
   wire _net_225;
   wire _net_221;
   wire _net_217;
   wire _net_215;
   wire _net_214;
   wire _net_213;
   wire _net_212;
   wire _net_211;
   wire _net_210;
   wire _net_209;
   wire _net_201;
   wire _net_193;
   wire _net_192;
   wire _net_191;
   wire _net_190;
   wire _net_189;
   wire _net_188;
   wire _net_184;
   wire _net_180;
   wire _net_178;
   wire _net_177;
   wire _net_176;
   wire _net_175;
   wire _net_174;
   wire _net_173;
   wire _net_172;
   wire _net_154;
   wire _net_129;
   wire _net_128;
   wire _net_127;
   wire _net_126;
   wire _net_125;
   wire _net_124;
   wire _net_123;
   wire _net_122;
   wire _net_121;
   wire _net_120;
   wire _net_119;
   wire _net_118;
   wire _net_117;
   wire _net_116;
   wire _net_115;
   wire _net_114;
   wire _net_113;

   // Assignments 

   // Module instantiations
   LOGIC1_X1 T0 (
	 );
   DFF_X1 L2199 (
	 );
   DFF_X1 L2198 (
	 );
   DFF_X1 L2197 (
	 );
   DFF_X1 L2196 (
	 );
   DFF_X1 L2195 (
	 );
   DFF_X1 L2194 (
	 );
   DFF_X1 L2193 (
	 );
   DFF_X1 L2192 (
	 );
   DFF_X1 L2191 (
	 );
   DFF_X1 L2190 (
	 );
   DFF_X1 L2189 (
	 );
   DFF_X1 L2188 (
	 );
   DFF_X1 L2187 (
	 );
   DFF_X1 L2186 (
	 );
   DFF_X1 L2185 (
	 );
   DFF_X1 L2184 (
	 );
   DFF_X1 L2183 (
	 );
   DFF_X1 L2182 (
	 );
   DFF_X1 L2181 (
	 );
   DFF_X1 L2180 (
	 );
   DFF_X1 L2179 (
	 );
   DFF_X1 L2178 (
	 );
   DFF_X1 L2177 (
	 );
   DFF_X1 L2176 (
	 );
   DFF_X1 L2175 (
	 );
   DFF_X1 L2174 (
	 );
   DFF_X1 L2173 (
	 );
   DFF_X1 L2172 (
	 );
   DFF_X1 L2171 (
	 );
   DFF_X1 L2170 (
	 );
   DFF_X1 L2169 (
	 );
   DFF_X1 L2168 (
	 );
   DFF_X1 L2167 (
	 );
   DFF_X1 L2166 (
	 );
   DFF_X1 L2165 (
	 );
   DFF_X1 L2164 (
	 );
   DFF_X1 L2163 (
	 );
   DFF_X1 L2162 (
	 );
   DFF_X1 L2161 (
	 );
   DFF_X1 L2160 (
	 );
   DFF_X1 L2159 (
	 );
   DFF_X1 L2158 (
	 );
   DFF_X1 L2157 (
	 );
   DFF_X1 L2156 (
	 );
   DFF_X1 L2155 (
	 );
   DFF_X1 L2154 (
	 );
   DFF_X1 L2153 (
	 );
   DFF_X1 L2152 (
	 );
   DFF_X1 L2151 (
	 );
   DFF_X1 L2150 (
	 );
   DFF_X1 L2149 (
	 );
   DFF_X1 L2148 (
	 );
   DFF_X1 L2147 (
	 );
   DFF_X1 L2146 (
	 );
   DFF_X1 L2145 (
	 );
   DFF_X1 L2144 (
	 );
   DFF_X1 L2143 (
	 );
   DFF_X1 L2142 (
	 );
   DFF_X1 L2141 (
	 );
   DFF_X1 L2140 (
	 );
   DFF_X1 L2139 (
	 );
   DFF_X1 L2138 (
	 );
   DFF_X1 L2137 (
	 );
   DFF_X1 L2136 (
	 );
   DFF_X1 L2135 (
	 );
   DFF_X1 L2134 (
	 );
   DFF_X1 L2133 (
	 );
   DFF_X1 L2132 (
	 );
   DFF_X1 L2131 (
	 );
   DFF_X1 L2130 (
	 );
   DFF_X1 L2129 (
	 );
   DFF_X1 L2128 (
	 );
   DFF_X1 L2127 (
	 );
   DFF_X1 L2126 (
	 );
   DFF_X1 L2125 (
	 );
   DFF_X1 L2124 (
	 );
   DFF_X1 L2123 (
	 );
   DFF_X1 L2122 (
	 );
   DFF_X1 L2121 (
	 );
   DFF_X1 L2120 (
	 );
   DFF_X1 L2119 (
	 );
   DFF_X1 L2118 (
	 );
   DFF_X1 L2117 (
	 );
   DFF_X1 L2116 (
	 );
   DFF_X1 L2115 (
	 );
   DFF_X1 L2114 (
	 );
   DFF_X1 L2113 (
	 );
   DFF_X1 L2112 (
	 );
   DFF_X1 L2111 (
	 );
   DFF_X1 L2110 (
	 );
   DFF_X1 L2109 (
	 );
   DFF_X1 L2108 (
	 );
   DFF_X1 L2107 (
	 );
   DFF_X1 L2106 (
	 );
   DFF_X1 L2105 (
	 );
   DFF_X1 L2104 (
	 );
   DFF_X1 L2103 (
	 );
   DFF_X1 L2102 (
	 );
   DFF_X1 L2101 (
	 );
   DFF_X1 L2100 (
	 );
   DFF_X1 L2099 (
	 );
   DFF_X1 L2098 (
	 );
   DFF_X1 L2097 (
	 );
   DFF_X1 L2096 (
	 );
   DFF_X1 L2095 (
	 );
   DFF_X1 L2094 (
	 );
   DFF_X1 L2093 (
	 );
   DFF_X1 L2092 (
	 );
   DFF_X1 L2091 (
	 );
   DFF_X1 L2090 (
	 );
   DFF_X1 L2089 (
	 );
   DFF_X1 L2088 (
	 );
   DFF_X1 L2087 (
	 );
   DFF_X1 L2086 (
	 );
   DFF_X1 L2085 (
	 );
   DFF_X1 L2084 (
	 );
   DFF_X1 L2083 (
	 );
   DFF_X1 L2082 (
	 );
   DFF_X1 L2081 (
	 );
   DFF_X1 L2080 (
	 );
   DFF_X1 L2079 (
	 );
   DFF_X1 L2078 (
	 );
   DFF_X1 L2077 (
	 );
   DFF_X1 L2076 (
	 );
   DFF_X1 L2075 (
	 );
   DFF_X1 L2074 (
	 );
   DFF_X1 L2073 (
	 );
   DFF_X1 L2072 (
	 );
   DFF_X1 L2071 (
	 );
   DFF_X1 L2070 (
	 );
   DFF_X1 L2069 (
	 );
   DFF_X1 L2068 (
	 );
   DFF_X1 L2067 (
	 );
   DFF_X1 L2066 (
	 );
   DFF_X1 L2065 (
	 );
   DFF_X1 L2064 (
	 );
   DFF_X1 L2063 (
	 );
   DFF_X1 L2062 (
	 );
   DFF_X1 L2061 (
	 );
   DFF_X1 L2060 (
	 );
   DFF_X1 L2059 (
	 );
   DFF_X1 L2058 (
	 );
   DFF_X1 L2057 (
	 );
   DFF_X1 L2056 (
	 );
   DFF_X1 L2055 (
	 );
   DFF_X1 L2054 (
	 );
   DFF_X1 L2053 (
	 );
   DFF_X1 L2052 (
	 );
   DFF_X1 L2051 (
	 );
   DFF_X1 L2050 (
	 );
   DFF_X1 L2049 (
	 );
   DFF_X1 L2048 (
	 );
   DFF_X1 L2047 (
	 );
   DFF_X1 L2046 (
	 );
   DFF_X1 L2045 (
	 );
   DFF_X1 L2044 (
	 );
   DFF_X1 L2043 (
	 );
   DFF_X1 L2042 (
	 );
   DFF_X1 L2041 (
	 );
   DFF_X1 L2040 (
	 );
   DFF_X1 L2039 (
	 );
   DFF_X1 L2038 (
	 );
   DFF_X1 L2037 (
	 );
   DFF_X1 L2036 (
	 );
   DFF_X1 L2035 (
	 );
   DFF_X1 L2034 (
	 );
   DFF_X1 L2033 (
	 );
   DFF_X1 L2032 (
	 );
   DFF_X1 L2031 (
	 );
   DFF_X1 L2030 (
	 );
   DFF_X1 L2029 (
	 );
   DFF_X1 L2028 (
	 );
   DFF_X1 L2027 (
	 );
   DFF_X1 L2026 (
	 );
   DFF_X1 L2025 (
	 );
   DFF_X1 L2024 (
	 );
   DFF_X1 L2023 (
	 );
   DFF_X1 L2022 (
	 );
   DFF_X1 L2021 (
	 );
   DFF_X1 L2020 (
	 );
   DFF_X1 L2019 (
	 );
   DFF_X1 L2018 (
	 );
   DFF_X1 L2017 (
	 );
   DFF_X1 L2016 (
	 );
   DFF_X1 L2015 (
	 );
   DFF_X1 L2014 (
	 );
   DFF_X1 L2013 (
	 );
   DFF_X1 L2012 (
	 );
   DFF_X1 L2011 (
	 );
   DFF_X1 L2010 (
	 );
   DFF_X1 L2009 (
	 );
   DFF_X1 L2008 (
	 );
   DFF_X1 L2007 (
	 );
   DFF_X1 L2006 (
	 );
   DFF_X1 L2005 (
	 );
   DFF_X1 L2004 (
	 );
   DFF_X1 L2003 (
	 );
   DFF_X1 L2002 (
	 );
   DFF_X1 L2001 (
	 );
   DFF_X1 L2000 (
	 );
   DFF_X1 L1999 (
	 );
   DFF_X1 L1998 (
	 );
   DFF_X1 L1997 (
	 );
   DFF_X1 L1996 (
	 );
   DFF_X1 L1995 (
	 );
   DFF_X1 L1994 (
	 );
   DFF_X1 L1993 (
	 );
   DFF_X1 L1992 (
	 );
   DFF_X1 L1991 (
	 );
   DFF_X1 L1990 (
	 );
   DFF_X1 L1989 (
	 );
   DFF_X1 L1988 (
	 );
   DFF_X1 L1987 (
	 );
   DFF_X1 L1986 (
	 );
   DFF_X1 L1985 (
	 );
   DFF_X1 L1984 (
	 );
   DFF_X1 L1983 (
	 );
   DFF_X1 L1982 (
	 );
   DFF_X1 L1981 (
	 );
   DFF_X1 L1980 (
	 );
   DFF_X1 L1979 (
	 );
   DFF_X1 L1978 (
	 );
   DFF_X1 L1977 (
	 );
   DFF_X1 L1976 (
	 );
   DFF_X1 L1975 (
	 );
   DFF_X1 L1974 (
	 );
   DFF_X1 L1973 (
	 );
   DFF_X1 L1972 (
	 );
   DFF_X1 L1971 (
	 );
   DFF_X1 L1970 (
	 );
   DFF_X1 L1969 (
	 );
   DFF_X1 L1968 (
	 );
   DFF_X1 L1967 (
	 );
   DFF_X1 L1966 (
	 );
   DFF_X1 L1965 (
	 );
   DFF_X1 L1964 (
	 );
   DFF_X1 L1963 (
	 );
   DFF_X1 L1962 (
	 );
   DFF_X1 L1961 (
	 );
   DFF_X1 L1960 (
	 );
   DFF_X1 L1959 (
	 );
   DFF_X1 L1958 (
	 );
   DFF_X1 L1957 (
	 );
   DFF_X1 L1956 (
	 );
   DFF_X1 L1955 (
	 );
   DFF_X1 L1954 (
	 );
   DFF_X1 L1953 (
	 );
   DFF_X1 L1952 (
	 );
   DFF_X1 L1951 (
	 );
   DFF_X1 L1950 (
	 );
   DFF_X1 L1949 (
	 );
   DFF_X1 L1948 (
	 );
   DFF_X1 L1947 (
	 );
   DFF_X1 L1946 (
	 );
   DFF_X1 L1945 (
	 );
   DFF_X1 L1944 (
	 );
   DFF_X1 L1943 (
	 );
   DFF_X1 L1942 (
	 );
   DFF_X1 L1941 (
	 );
   DFF_X1 L1940 (
	 );
   DFF_X1 L1939 (
	 );
   DFF_X1 L1938 (
	 );
   DFF_X1 L1937 (
	 );
   DFF_X1 L1936 (
	 );
   DFF_X1 L1935 (
	 );
   DFF_X1 L1934 (
	 );
   DFF_X1 L1933 (
	 );
   DFF_X1 L1932 (
	 );
   DFF_X1 L1931 (
	 );
   DFF_X1 L1930 (
	 );
   DFF_X1 L1929 (
	 );
   DFF_X1 L1928 (
	 );
   DFF_X1 L1927 (
	 );
   DFF_X1 L1926 (
	 );
   DFF_X1 L1925 (
	 );
   DFF_X1 L1924 (
	 );
   DFF_X1 L1923 (
	 );
   DFF_X1 L1922 (
	 );
   DFF_X1 L1921 (
	 );
   DFF_X1 L1920 (
	 );
   DFF_X1 L1919 (
	 );
   DFF_X1 L1918 (
	 );
   DFF_X1 L1917 (
	 );
   DFF_X1 L1916 (
	 );
   DFF_X1 L1915 (
	 );
   DFF_X1 L1914 (
	 );
   DFF_X1 L1913 (
	 );
   DFF_X1 L1912 (
	 );
   DFF_X1 L1911 (
	 );
   DFF_X1 L1910 (
	 );
   DFF_X1 L1909 (
	 );
   DFF_X1 L1908 (
	 );
   DFF_X1 L1907 (
	 );
   DFF_X1 L1906 (
	 );
   DFF_X1 L1905 (
	 );
   DFF_X1 L1904 (
	 );
   DFF_X1 L1903 (
	 );
   DFF_X1 L1902 (
	 );
   DFF_X1 L1901 (
	 );
   DFF_X1 L1900 (
	 );
   DFF_X1 L1899 (
	 );
   DFF_X1 L1898 (
	 );
   DFF_X1 L1897 (
	 );
   DFF_X1 L1896 (
	 );
   DFF_X1 L1895 (
	 );
   DFF_X1 L1894 (
	 );
   DFF_X1 L1893 (
	 );
   DFF_X1 L1892 (
	 );
   DFF_X1 L1891 (
	 );
   DFF_X1 L1890 (
	 );
   DFF_X1 L1889 (
	 );
   DFF_X1 L1888 (
	 );
   DFF_X1 L1887 (
	 );
   DFF_X1 L1886 (
	 );
   DFF_X1 L1885 (
	 );
   DFF_X1 L1884 (
	 );
   DFF_X1 L1883 (
	 );
   DFF_X1 L1882 (
	 );
   DFF_X1 L1881 (
	 );
   DFF_X1 L1880 (
	 );
   DFF_X1 L1879 (
	 );
   DFF_X1 L1878 (
	 );
   DFF_X1 L1877 (
	 );
   DFF_X1 L1876 (
	 );
   DFF_X1 L1875 (
	 );
   DFF_X1 L1874 (
	 );
   DFF_X1 L1873 (
	 );
   DFF_X1 L1872 (
	 );
   DFF_X1 L1871 (
	 );
   DFF_X1 L1870 (
	 );
   DFF_X1 L1869 (
	 );
   DFF_X1 L1868 (
	 );
   DFF_X1 L1867 (
	 );
   DFF_X1 L1866 (
	 );
   DFF_X1 L1865 (
	 );
   DFF_X1 L1864 (
	 );
   DFF_X1 L1863 (
	 );
   DFF_X1 L1862 (
	 );
   DFF_X1 L1861 (
	 );
   DFF_X1 L1860 (
	 );
   DFF_X1 L1859 (
	 );
   DFF_X1 L1858 (
	 );
   DFF_X1 L1857 (
	 );
   DFF_X1 L1856 (
	 );
   DFF_X1 L1855 (
	 );
   DFF_X1 L1854 (
	 );
   DFF_X1 L1853 (
	 );
   DFF_X1 L1852 (
	 );
   DFF_X1 L1851 (
	 );
   DFF_X1 L1850 (
	 );
   DFF_X1 L1849 (
	 );
   DFF_X1 L1848 (
	 );
   DFF_X1 L1847 (
	 );
   DFF_X1 L1846 (
	 );
   DFF_X1 L1845 (
	 );
   DFF_X1 L1844 (
	 );
   DFF_X1 L1843 (
	 );
   DFF_X1 L1842 (
	 );
   DFF_X1 L1841 (
	 );
   DFF_X1 L1840 (
	 );
   DFF_X1 L1839 (
	 );
   DFF_X1 L1838 (
	 );
   DFF_X1 L1837 (
	 );
   DFF_X1 L1836 (
	 );
   DFF_X1 L1835 (
	 );
   DFF_X1 L1834 (
	 );
   DFF_X1 L1833 (
	 );
   DFF_X1 L1832 (
	 );
   DFF_X1 L1831 (
	 );
   DFF_X1 L1830 (
	 );
   DFF_X1 L1829 (
	 );
   DFF_X1 L1828 (
	 );
   DFF_X1 L1827 (
	 );
   DFF_X1 L1826 (
	 );
   DFF_X1 L1825 (
	 );
   DFF_X1 L1824 (
	 );
   DFF_X1 L1823 (
	 );
   DFF_X1 L1822 (
	 );
   DFF_X1 L1821 (
	 );
   DFF_X1 L1820 (
	 );
   DFF_X1 L1819 (
	 );
   DFF_X1 L1818 (
	 );
   DFF_X1 L1817 (
	 );
   DFF_X1 L1816 (
	 );
   DFF_X1 L1815 (
	 );
   DFF_X1 L1814 (
	 );
   DFF_X1 L1813 (
	 );
   DFF_X1 L1812 (
	 );
   DFF_X1 L1811 (
	 );
   DFF_X1 L1810 (
	 );
   DFF_X1 L1809 (
	 );
   DFF_X1 L1808 (
	 );
   DFF_X1 L1807 (
	 );
   DFF_X1 L1806 (
	 );
   DFF_X1 L1805 (
	 );
   DFF_X1 L1804 (
	 );
   DFF_X1 L1803 (
	 );
   DFF_X1 L1802 (
	 );
   DFF_X1 L1801 (
	 );
   DFF_X1 L1800 (
	 );
   DFF_X1 L1799 (
	 );
   DFF_X1 L1798 (
	 );
   DFF_X1 L1797 (
	 );
   DFF_X1 L1796 (
	 );
   DFF_X1 L1795 (
	 );
   DFF_X1 L1794 (
	 );
   DFF_X1 L1793 (
	 );
   DFF_X1 L1792 (
	 );
   DFF_X1 L1791 (
	 );
   DFF_X1 L1790 (
	 );
   DFF_X1 L1789 (
	 );
   DFF_X1 L1788 (
	 );
   DFF_X1 L1787 (
	 );
   DFF_X1 L1786 (
	 );
   DFF_X1 L1785 (
	 );
   DFF_X1 L1784 (
	 );
   DFF_X1 L1783 (
	 );
   DFF_X1 L1782 (
	 );
   DFF_X1 L1781 (
	 );
   DFF_X1 L1780 (
	 );
   DFF_X1 L1779 (
	 );
   DFF_X1 L1778 (
	 );
   DFF_X1 L1777 (
	 );
   DFF_X1 L1776 (
	 );
   DFF_X1 L1775 (
	 );
   DFF_X1 L1774 (
	 );
   DFF_X1 L1773 (
	 );
   DFF_X1 L1772 (
	 );
   DFF_X1 L1771 (
	 );
   DFF_X1 L1770 (
	 );
   DFF_X1 L1769 (
	 );
   DFF_X1 L1768 (
	 );
   DFF_X1 L1767 (
	 );
   DFF_X1 L1766 (
	 );
   DFF_X1 L1765 (
	 );
   DFF_X1 L1764 (
	 );
   DFF_X1 L1763 (
	 );
   DFF_X1 L1762 (
	 );
   DFF_X1 L1761 (
	 );
   DFF_X1 L1760 (
	 );
   DFF_X1 L1759 (
	 );
   DFF_X1 L1758 (
	 );
   DFF_X1 L1757 (
	 );
   DFF_X1 L1756 (
	 );
   DFF_X1 L1755 (
	 );
   DFF_X1 L1754 (
	 );
   DFF_X1 L1753 (
	 );
   DFF_X1 L1752 (
	 );
   DFF_X1 L1751 (
	 );
   DFF_X1 L1750 (
	 );
   DFF_X1 L1749 (
	 );
   DFF_X1 L1748 (
	 );
   DFF_X1 L1747 (
	 );
   DFF_X1 L1746 (
	 );
   DFF_X1 L1745 (
	 );
   DFF_X1 L1744 (
	 );
   DFF_X1 L1743 (
	 );
   DFF_X1 L1742 (
	 );
   DFF_X1 L1741 (
	 );
   DFF_X1 L1740 (
	 );
   DFF_X1 L1739 (
	 );
   DFF_X1 L1738 (
	 );
   DFF_X1 L1737 (
	 );
   DFF_X1 L1736 (
	 );
   DFF_X1 L1735 (
	 );
   DFF_X1 L1734 (
	 );
   DFF_X1 L1733 (
	 );
   DFF_X1 L1732 (
	 );
   DFF_X1 L1731 (
	 );
   DFF_X1 L1730 (
	 );
   DFF_X1 L1729 (
	 );
   DFF_X1 L1728 (
	 );
   DFF_X1 L1727 (
	 );
   DFF_X1 L1726 (
	 );
   DFF_X1 L1725 (
	 );
   DFF_X1 L1724 (
	 );
   DFF_X1 L1723 (
	 );
   DFF_X1 L1722 (
	 );
   DFF_X1 L1721 (
	 );
   DFF_X1 L1720 (
	 );
   DFF_X1 L1719 (
	 );
   DFF_X1 L1718 (
	 );
   DFF_X1 L1717 (
	 );
   DFF_X1 L1716 (
	 );
   DFF_X1 L1715 (
	 );
   DFF_X1 L1714 (
	 );
   DFF_X1 L1713 (
	 );
   DFF_X1 L1712 (
	 );
   DFF_X1 L1711 (
	 );
   DFF_X1 L1710 (
	 );
   DFF_X1 L1709 (
	 );
   DFF_X1 L1708 (
	 );
   DFF_X1 L1707 (
	 );
   DFF_X1 L1706 (
	 );
   DFF_X1 L1705 (
	 );
   DFF_X1 L1704 (
	 );
   DFF_X1 L1703 (
	 );
   DFF_X1 L1702 (
	 );
   DFF_X1 L1701 (
	 );
   DFF_X1 L1700 (
	 );
   DFF_X1 L1699 (
	 );
   DFF_X1 L1698 (
	 );
   DFF_X1 L1697 (
	 );
   DFF_X1 L1696 (
	 );
   DFF_X1 L1695 (
	 );
   DFF_X1 L1694 (
	 );
   DFF_X1 L1693 (
	 );
   DFF_X1 L1692 (
	 );
   DFF_X1 L1691 (
	 );
   DFF_X1 L1690 (
	 );
   DFF_X1 L1689 (
	 );
   DFF_X1 L1688 (
	 );
   DFF_X1 L1687 (
	 );
   DFF_X1 L1686 (
	 );
   DFF_X1 L1685 (
	 );
   DFF_X1 L1684 (
	 );
   DFF_X1 L1683 (
	 );
   DFF_X1 L1682 (
	 );
   DFF_X1 L1681 (
	 );
   DFF_X1 L1680 (
	 );
   DFF_X1 L1679 (
	 );
   DFF_X1 L1678 (
	 );
   DFF_X1 L1677 (
	 );
   DFF_X1 L1676 (
	 );
   DFF_X1 L1675 (
	 );
   DFF_X1 L1674 (
	 );
   DFF_X1 L1673 (
	 );
   DFF_X1 L1672 (
	 );
   DFF_X1 L1671 (
	 );
   DFF_X1 L1670 (
	 );
   DFF_X1 L1669 (
	 );
   DFF_X1 L1668 (
	 );
   DFF_X1 L1667 (
	 );
   DFF_X1 L1666 (
	 );
   DFF_X1 L1665 (
	 );
   DFF_X1 L1664 (
	 );
   DFF_X1 L1663 (
	 );
   DFF_X1 L1662 (
	 );
   DFF_X1 L1661 (
	 );
   DFF_X1 L1660 (
	 );
   DFF_X1 L1659 (
	 );
   DFF_X1 L1658 (
	 );
   DFF_X1 L1657 (
	 );
   DFF_X1 L1656 (
	 );
   DFF_X1 L1655 (
	 );
   DFF_X1 L1654 (
	 );
   DFF_X1 L1653 (
	 );
   DFF_X1 L1652 (
	 );
   DFF_X1 L1651 (
	 );
   DFF_X1 L1650 (
	 );
   DFF_X1 L1649 (
	 );
   DFF_X1 L1648 (
	 );
   DFF_X1 L1647 (
	 );
   DFF_X1 L1646 (
	 );
   DFF_X1 L1645 (
	 );
   DFF_X1 L1644 (
	 );
   DFF_X1 L1643 (
	 );
   DFF_X1 L1642 (
	 );
   DFF_X1 L1641 (
	 );
   DFF_X1 L1640 (
	 );
   DFF_X1 L1639 (
	 );
   DFF_X1 L1638 (
	 );
   DFF_X1 L1637 (
	 );
   DFF_X1 L1636 (
	 );
   DFF_X1 L1635 (
	 );
   DFF_X1 L1634 (
	 );
   DFF_X1 L1633 (
	 );
   DFF_X1 L1632 (
	 );
   DFF_X1 L1631 (
	 );
   DFF_X1 L1630 (
	 );
   DFF_X1 L1629 (
	 );
   DFF_X1 L1628 (
	 );
   DFF_X1 L1627 (
	 );
   DFF_X1 L1626 (
	 );
   DFF_X1 L1625 (
	 );
   DFF_X1 L1624 (
	 );
   DFF_X1 L1623 (
	 );
   DFF_X1 L1622 (
	 );
   DFF_X1 L1621 (
	 );
   DFF_X1 L1620 (
	 );
   DFF_X1 L1619 (
	 );
   DFF_X1 L1618 (
	 );
   DFF_X1 L1617 (
	 );
   DFF_X1 L1616 (
	 );
   DFF_X1 L1615 (
	 );
   DFF_X1 L1614 (
	 );
   DFF_X1 L1613 (
	 );
   DFF_X1 L1612 (
	 );
   DFF_X1 L1611 (
	 );
   DFF_X1 L1610 (
	 );
   DFF_X1 L1609 (
	 );
   DFF_X1 L1608 (
	 );
   DFF_X1 L1607 (
	 );
   DFF_X1 L1606 (
	 );
   DFF_X1 L1605 (
	 );
   DFF_X1 L1604 (
	 );
   DFF_X1 L1603 (
	 );
   DFF_X1 L1602 (
	 );
   DFF_X1 L1601 (
	 );
   DFF_X1 L1600 (
	 );
   DFF_X1 L1599 (
	 );
   DFF_X1 L1598 (
	 );
   DFF_X1 L1597 (
	 );
   DFF_X1 L1596 (
	 );
   DFF_X1 L1595 (
	 );
   DFF_X1 L1594 (
	 );
   DFF_X1 L1593 (
	 );
   DFF_X1 L1592 (
	 );
   DFF_X1 L1591 (
	 );
   DFF_X1 L1590 (
	 );
   DFF_X1 L1589 (
	 );
   DFF_X1 L1588 (
	 );
   DFF_X1 L1587 (
	 );
   DFF_X1 L1586 (
	 );
   DFF_X1 L1585 (
	 );
   DFF_X1 L1584 (
	 );
   DFF_X1 L1583 (
	 );
   DFF_X1 L1582 (
	 );
   DFF_X1 L1581 (
	 );
   DFF_X1 L1580 (
	 );
   DFF_X1 L1579 (
	 );
   DFF_X1 L1578 (
	 );
   DFF_X1 L1577 (
	 );
   DFF_X1 L1576 (
	 );
   DFF_X1 L1575 (
	 );
   DFF_X1 L1574 (
	 );
   DFF_X1 L1573 (
	 );
   DFF_X1 L1572 (
	 );
   DFF_X1 L1571 (
	 );
   DFF_X1 L1570 (
	 );
   DFF_X1 L1569 (
	 );
   DFF_X1 L1568 (
	 );
   DFF_X1 L1567 (
	 );
   DFF_X1 L1566 (
	 );
   DFF_X1 L1565 (
	 );
   DFF_X1 L1564 (
	 );
   DFF_X1 L1563 (
	 );
   DFF_X1 L1562 (
	 );
   DFF_X1 L1561 (
	 );
   DFF_X1 L1560 (
	 );
   DFF_X1 L1559 (
	 );
   DFF_X1 L1558 (
	 );
   DFF_X1 L1557 (
	 );
   DFF_X1 L1556 (
	 );
   DFF_X1 L1555 (
	 );
   DFF_X1 L1554 (
	 );
   DFF_X1 L1553 (
	 );
   DFF_X1 L1552 (
	 );
   DFF_X1 L1551 (
	 );
   DFF_X1 L1550 (
	 );
   DFF_X1 L1549 (
	 );
   DFF_X1 L1548 (
	 );
   DFF_X1 L1547 (
	 );
   DFF_X1 L1546 (
	 );
   DFF_X1 L1545 (
	 );
   DFF_X1 L1544 (
	 );
   DFF_X1 L1543 (
	 );
   DFF_X1 L1542 (
	 );
   DFF_X1 L1541 (
	 );
   DFF_X1 L1540 (
	 );
   DFF_X1 L1539 (
	 );
   DFF_X1 L1538 (
	 );
   DFF_X1 L1537 (
	 );
   DFF_X1 L1536 (
	 );
   DFF_X1 L1535 (
	 );
   DFF_X1 L1534 (
	 );
   DFF_X1 L1533 (
	 );
   DFF_X1 L1532 (
	 );
   DFF_X1 L1531 (
	 );
   DFF_X1 L1530 (
	 );
   DFF_X1 L1529 (
	 );
   DFF_X1 L1528 (
	 );
   DFF_X1 L1527 (
	 );
   DFF_X1 L1526 (
	 );
   DFF_X1 L1525 (
	 );
   DFF_X1 L1524 (
	 );
   DFF_X1 L1523 (
	 );
   DFF_X1 L1522 (
	 );
   DFF_X1 L1521 (
	 );
   DFF_X1 L1520 (
	 );
   DFF_X1 L1519 (
	 );
   DFF_X1 L1518 (
	 );
   DFF_X1 L1517 (
	 );
   DFF_X1 L1516 (
	 );
   DFF_X1 L1515 (
	 );
   DFF_X1 L1514 (
	 );
   DFF_X1 L1513 (
	 );
   DFF_X1 L1512 (
	 );
   DFF_X1 L1511 (
	 );
   DFF_X1 L1510 (
	 );
   DFF_X1 L1509 (
	 );
   DFF_X1 L1508 (
	 );
   DFF_X1 L1507 (
	 );
   DFF_X1 L1506 (
	 );
   DFF_X1 L1505 (
	 );
   DFF_X1 L1504 (
	 );
   DFF_X1 L1503 (
	 );
   DFF_X1 L1502 (
	 );
   DFF_X1 L1501 (
	 );
   DFF_X1 L1500 (
	 );
   DFF_X1 L1499 (
	 );
   DFF_X1 L1498 (
	 );
   DFF_X1 L1497 (
	 );
   DFF_X1 L1496 (
	 );
   DFF_X1 L1495 (
	 );
   DFF_X1 L1494 (
	 );
   DFF_X1 L1493 (
	 );
   DFF_X1 L1492 (
	 );
   DFF_X1 L1491 (
	 );
   DFF_X1 L1490 (
	 );
   DFF_X1 L1489 (
	 );
   DFF_X1 L1488 (
	 );
   DFF_X1 L1487 (
	 );
   DFF_X1 L1486 (
	 );
   DFF_X1 L1485 (
	 );
   DFF_X1 L1484 (
	 );
   DFF_X1 L1483 (
	 );
   DFF_X1 L1482 (
	 );
   DFF_X1 L1481 (
	 );
   DFF_X1 L1480 (
	 );
   DFF_X1 L1479 (
	 );
   DFF_X1 L1478 (
	 );
   DFF_X1 L1477 (
	 );
   DFF_X1 L1476 (
	 );
   DFF_X1 L1475 (
	 );
   DFF_X1 L1474 (
	 );
   DFF_X1 L1473 (
	 );
   DFF_X1 L1472 (
	 );
   DFF_X1 L1471 (
	 );
   DFF_X1 L1470 (
	 );
   DFF_X1 L1469 (
	 );
   DFF_X1 L1468 (
	 );
   DFF_X1 L1467 (
	 );
   DFF_X1 L1466 (
	 );
   DFF_X1 L1465 (
	 );
   DFF_X1 L1464 (
	 );
   DFF_X1 L1463 (
	 );
   DFF_X1 L1462 (
	 );
   DFF_X1 L1461 (
	 );
   DFF_X1 L1460 (
	 );
   DFF_X1 L1459 (
	 );
   DFF_X1 L1458 (
	 );
   DFF_X1 L1457 (
	 );
   DFF_X1 L1456 (
	 );
   DFF_X1 L1455 (
	 );
   DFF_X1 L1454 (
	 );
   DFF_X1 L1453 (
	 );
   DFF_X1 L1452 (
	 );
   DFF_X1 L1451 (
	 );
   DFF_X1 L1450 (
	 );
   DFF_X1 L1449 (
	 );
   DFF_X1 L1448 (
	 );
   DFF_X1 L1447 (
	 );
   DFF_X1 L1446 (
	 );
   DFF_X1 L1445 (
	 );
   DFF_X1 L1444 (
	 );
   DFF_X1 L1443 (
	 );
   DFF_X1 L1442 (
	 );
   DFF_X1 L1441 (
	 );
   DFF_X1 L1440 (
	 );
   DFF_X1 L1439 (
	 );
   DFF_X1 L1438 (
	 );
   DFF_X1 L1437 (
	 );
   DFF_X1 L1436 (
	 );
   DFF_X1 L1435 (
	 );
   DFF_X1 L1434 (
	 );
   DFF_X1 L1433 (
	 );
   DFF_X1 L1432 (
	 );
   DFF_X1 L1431 (
	 );
   DFF_X1 L1430 (
	 );
   DFF_X1 L1429 (
	 );
   DFF_X1 L1428 (
	 );
   DFF_X1 L1427 (
	 );
   DFF_X1 L1426 (
	 );
   DFF_X1 L1425 (
	 );
   DFF_X1 L1424 (
	 );
   DFF_X1 L1423 (
	 );
   DFF_X1 L1422 (
	 );
   DFF_X1 L1421 (
	 );
   DFF_X1 L1420 (
	 );
   DFF_X1 L1419 (
	 );
   DFF_X1 L1418 (
	 );
   DFF_X1 L1417 (
	 );
   DFF_X1 L1416 (
	 );
   DFF_X1 L1415 (
	 );
   DFF_X1 L1414 (
	 );
   DFF_X1 L1413 (
	 );
   DFF_X1 L1412 (
	 );
   DFF_X1 L1411 (
	 );
   DFF_X1 L1410 (
	 );
   DFF_X1 L1409 (
	 );
   DFF_X1 L1408 (
	 );
   DFF_X1 L1407 (
	 );
   DFF_X1 L1406 (
	 );
   DFF_X1 L1405 (
	 );
   DFF_X1 L1404 (
	 );
   DFF_X1 L1403 (
	 );
   DFF_X1 L1402 (
	 );
   DFF_X1 L1401 (
	 );
   DFF_X1 L1400 (
	 );
   DFF_X1 L1399 (
	 );
   DFF_X1 L1398 (
	 );
   DFF_X1 L1397 (
	 );
   DFF_X1 L1396 (
	 );
   DFF_X1 L1395 (
	 );
   DFF_X1 L1394 (
	 );
   DFF_X1 L1393 (
	 );
   DFF_X1 L1392 (
	 );
   DFF_X1 L1391 (
	 );
   DFF_X1 L1390 (
	 );
   DFF_X1 L1389 (
	 );
   DFF_X1 L1388 (
	 );
   DFF_X1 L1387 (
	 );
   DFF_X1 L1386 (
	 );
   DFF_X1 L1385 (
	 );
   DFF_X1 L1384 (
	 );
   DFF_X1 L1383 (
	 );
   DFF_X1 L1382 (
	 );
   DFF_X1 L1381 (
	 );
   DFF_X1 L1380 (
	 );
   DFF_X1 L1379 (
	 );
   DFF_X1 L1378 (
	 );
   DFF_X1 L1377 (
	 );
   DFF_X1 L1376 (
	 );
   DFF_X1 L1375 (
	 );
   DFF_X1 L1374 (
	 );
   DFF_X1 L1373 (
	 );
   DFF_X1 L1372 (
	 );
   DFF_X1 L1371 (
	 );
   DFF_X1 L1370 (
	 );
   DFF_X1 L1369 (
	 );
   DFF_X1 L1368 (
	 );
   DFF_X1 L1367 (
	 );
   DFF_X1 L1366 (
	 );
   DFF_X1 L1365 (
	 );
   DFF_X1 L1364 (
	 );
   DFF_X1 L1363 (
	 );
   DFF_X1 L1362 (
	 );
   DFF_X1 L1361 (
	 );
   DFF_X1 L1360 (
	 );
   DFF_X1 L1359 (
	 );
   DFF_X1 L1358 (
	 );
   DFF_X1 L1357 (
	 );
   DFF_X1 L1356 (
	 );
   DFF_X1 L1355 (
	 );
   DFF_X1 L1354 (
	 );
   DFF_X1 L1353 (
	 );
   DFF_X1 L1352 (
	 );
   DFF_X1 L1351 (
	 );
   DFF_X1 L1350 (
	 );
   DFF_X1 L1349 (
	 );
   DFF_X1 L1348 (
	 );
   DFF_X1 L1347 (
	 );
   DFF_X1 L1346 (
	 );
   DFF_X1 L1345 (
	 );
   DFF_X1 L1344 (
	 );
   DFF_X1 L1343 (
	 );
   DFF_X1 L1342 (
	 );
   DFF_X1 L1341 (
	 );
   DFF_X1 L1340 (
	 );
   DFF_X1 L1339 (
	 );
   DFF_X1 L1338 (
	 );
   DFF_X1 L1337 (
	 );
   DFF_X1 L1336 (
	 );
   DFF_X1 L1335 (
	 );
   DFF_X1 L1334 (
	 );
   DFF_X1 L1333 (
	 );
   DFF_X1 L1332 (
	 );
   DFF_X1 L1331 (
	 );
   DFF_X1 L1330 (
	 );
   DFF_X1 L1329 (
	 );
   DFF_X1 L1328 (
	 );
   DFF_X1 L1327 (
	 );
   DFF_X1 L1326 (
	 );
   DFF_X1 L1325 (
	 );
   DFF_X1 L1324 (
	 );
   DFF_X1 L1323 (
	 );
   DFF_X1 L1322 (
	 );
   DFF_X1 L1321 (
	 );
   DFF_X1 L1320 (
	 );
   DFF_X1 L1319 (
	 );
   DFF_X1 L1318 (
	 );
   DFF_X1 L1317 (
	 );
   DFF_X1 L1316 (
	 );
   DFF_X1 L1315 (
	 );
   DFF_X1 L1314 (
	 );
   DFF_X1 L1313 (
	 );
   DFF_X1 L1312 (
	 );
   DFF_X1 L1311 (
	 );
   DFF_X1 L1310 (
	 );
   DFF_X1 L1309 (
	 );
   DFF_X1 L1308 (
	 );
   DFF_X1 L1307 (
	 );
   DFF_X1 L1306 (
	 );
   DFF_X1 L1305 (
	 );
   DFF_X1 L1304 (
	 );
   DFF_X1 L1303 (
	 );
   DFF_X1 L1302 (
	 );
   DFF_X1 L1301 (
	 );
   DFF_X1 L1300 (
	 );
   DFF_X1 L1299 (
	 );
   DFF_X1 L1298 (
	 );
   DFF_X1 L1297 (
	 );
   DFF_X1 L1296 (
	 );
   DFF_X1 L1295 (
	 );
   DFF_X1 L1294 (
	 );
   DFF_X1 L1293 (
	 );
   DFF_X1 L1292 (
	 );
   DFF_X1 L1291 (
	 );
   DFF_X1 L1290 (
	 );
   DFF_X1 L1289 (
	 );
   DFF_X1 L1288 (
	 );
   DFF_X1 L1287 (
	 );
   DFF_X1 L1286 (
	 );
   DFF_X1 L1285 (
	 );
   DFF_X1 L1284 (
	 );
   DFF_X1 L1283 (
	 );
   DFF_X1 L1282 (
	 );
   DFF_X1 L1281 (
	 );
   DFF_X1 L1280 (
	 );
   DFF_X1 L1279 (
	 );
   DFF_X1 L1278 (
	 );
   DFF_X1 L1277 (
	 );
   DFF_X1 L1276 (
	 );
   DFF_X1 L1275 (
	 );
   DFF_X1 L1274 (
	 );
   DFF_X1 L1273 (
	 );
   DFF_X1 L1272 (
	 );
   DFF_X1 L1271 (
	 );
   DFF_X1 L1270 (
	 );
   DFF_X1 L1269 (
	 );
   DFF_X1 L1268 (
	 );
   DFF_X1 L1267 (
	 );
   DFF_X1 L1266 (
	 );
   DFF_X1 L1265 (
	 );
   DFF_X1 L1264 (
	 );
   DFF_X1 L1263 (
	 );
   DFF_X1 L1262 (
	 );
   DFF_X1 L1261 (
	 );
   DFF_X1 L1260 (
	 );
   DFF_X1 L1259 (
	 );
   DFF_X1 L1258 (
	 );
   DFF_X1 L1257 (
	 );
   DFF_X1 L1256 (
	 );
   DFF_X1 L1255 (
	 );
   DFF_X1 L1254 (
	 );
   DFF_X1 L1253 (
	 );
   DFF_X1 L1252 (
	 );
   DFF_X1 L1251 (
	 );
   DFF_X1 L1250 (
	 );
   DFF_X1 L1249 (
	 );
   DFF_X1 L1248 (
	 );
   DFF_X1 L1247 (
	 );
   DFF_X1 L1246 (
	 );
   DFF_X1 L1245 (
	 );
   DFF_X1 L1244 (
	 );
   DFF_X1 L1243 (
	 );
   DFF_X1 L1242 (
	 );
   DFF_X1 L1241 (
	 );
   DFF_X1 L1240 (
	 );
   DFF_X1 L1239 (
	 );
   DFF_X1 L1238 (
	 );
   DFF_X1 L1237 (
	 );
   DFF_X1 L1236 (
	 );
   DFF_X1 L1235 (
	 );
   DFF_X1 L1234 (
	 );
   DFF_X1 L1233 (
	 );
   DFF_X1 L1232 (
	 );
   DFF_X1 L1231 (
	 );
   DFF_X1 L1230 (
	 );
   DFF_X1 L1229 (
	 );
   DFF_X1 L1228 (
	 );
   DFF_X1 L1227 (
	 );
   DFF_X1 L1226 (
	 );
   DFF_X1 L1225 (
	 );
   DFF_X1 L1224 (
	 );
   DFF_X1 L1223 (
	 );
   DFF_X1 L1222 (
	 );
   DFF_X1 L1221 (
	 );
   DFF_X1 L1220 (
	 );
   DFF_X1 L1219 (
	 );
   DFF_X1 L1218 (
	 );
   DFF_X1 L1217 (
	 );
   DFF_X1 L1216 (
	 );
   DFF_X1 L1215 (
	 );
   DFF_X1 L1214 (
	 );
   DFF_X1 L1213 (
	 );
   DFF_X1 L1212 (
	 );
   DFF_X1 L1211 (
	 );
   DFF_X1 L1210 (
	 );
   DFF_X1 L1209 (
	 );
   DFF_X1 L1208 (
	 );
   DFF_X1 L1207 (
	 );
   DFF_X1 L1206 (
	 );
   DFF_X1 L1205 (
	 );
   DFF_X1 L1204 (
	 );
   DFF_X1 L1203 (
	 );
   DFF_X1 L1202 (
	 );
   DFF_X1 L1201 (
	 );
   DFF_X1 L1200 (
	 );
   DFF_X1 L1199 (
	 );
   DFF_X1 L1198 (
	 );
   DFF_X1 L1197 (
	 );
   DFF_X1 L1196 (
	 );
   DFF_X1 L1195 (
	 );
   DFF_X1 L1194 (
	 );
   DFF_X1 L1193 (
	 );
   DFF_X1 L1192 (
	 );
   DFF_X1 L1191 (
	 );
   DFF_X1 L1190 (
	 );
   DFF_X1 L1189 (
	 );
   DFF_X1 L1188 (
	 );
   DFF_X1 L1187 (
	 );
   DFF_X1 L1186 (
	 );
   DFF_X1 L1185 (
	 );
   DFF_X1 L1184 (
	 );
   DFF_X1 L1183 (
	 );
   DFF_X1 L1182 (
	 );
   DFF_X1 L1181 (
	 );
   DFF_X1 L1180 (
	 );
   DFF_X1 L1179 (
	 );
   DFF_X1 L1178 (
	 );
   DFF_X1 L1177 (
	 );
   DFF_X1 L1176 (
	 );
   DFF_X1 L1175 (
	 );
   DFF_X1 L1174 (
	 );
   DFF_X1 L1173 (
	 );
   DFF_X1 L1172 (
	 );
   DFF_X1 L1171 (
	 );
   DFF_X1 L1170 (
	 );
   DFF_X1 L1169 (
	 );
   DFF_X1 L1168 (
	 );
   DFF_X1 L1167 (
	 );
   DFF_X1 L1166 (
	 );
   DFF_X1 L1165 (
	 );
   DFF_X1 L1164 (
	 );
   DFF_X1 L1163 (
	 );
   DFF_X1 L1162 (
	 );
   DFF_X1 L1161 (
	 );
   DFF_X1 L1160 (
	 );
   DFF_X1 L1159 (
	 );
   DFF_X1 L1158 (
	 );
   DFF_X1 L1157 (
	 );
   DFF_X1 L1156 (
	 );
   DFF_X1 L1155 (
	 );
   DFF_X1 L1154 (
	 );
   DFF_X1 L1153 (
	 );
   DFF_X1 L1152 (
	 );
   DFF_X1 L1151 (
	 );
   DFF_X1 L1150 (
	 );
   DFF_X1 L1149 (
	 );
   DFF_X1 L1148 (
	 );
   DFF_X1 L1147 (
	 );
   DFF_X1 L1146 (
	 );
   DFF_X1 L1145 (
	 );
   DFF_X1 L1144 (
	 );
   DFF_X1 L1143 (
	 );
   DFF_X1 L1142 (
	 );
   DFF_X1 L1141 (
	 );
   DFF_X1 L1140 (
	 );
   DFF_X1 L1139 (
	 );
   DFF_X1 L1138 (
	 );
   DFF_X1 L1137 (
	 );
   DFF_X1 L1136 (
	 );
   DFF_X1 L1135 (
	 );
   DFF_X1 L1134 (
	 );
   DFF_X1 L1133 (
	 );
   DFF_X1 L1132 (
	 );
   DFF_X1 L1131 (
	 );
   DFF_X1 L1130 (
	 );
   DFF_X1 L1129 (
	 );
   DFF_X1 L1128 (
	 );
   DFF_X1 L1127 (
	 );
   DFF_X1 L1126 (
	 );
   DFF_X1 L1125 (
	 );
   DFF_X1 L1124 (
	 );
   DFF_X1 L1123 (
	 );
   DFF_X1 L1122 (
	 );
   DFF_X1 L1121 (
	 );
   DFF_X1 L1120 (
	 );
   DFF_X1 L1119 (
	 );
   DFF_X1 L1118 (
	 );
   DFF_X1 L1117 (
	 );
   DFF_X1 L1116 (
	 );
   DFF_X1 L1115 (
	 );
   DFF_X1 L1114 (
	 );
   DFF_X1 L1113 (
	 );
   DFF_X1 L1112 (
	 );
   DFF_X1 L1111 (
	 );
   DFF_X1 L1110 (
	 );
   DFF_X1 L1109 (
	 );
   DFF_X1 L1108 (
	 );
   DFF_X1 L1107 (
	 );
   DFF_X1 L1106 (
	 );
   DFF_X1 L1105 (
	 );
   DFF_X1 L1104 (
	 );
   DFF_X1 L1103 (
	 );
   DFF_X1 L1102 (
	 );
   DFF_X1 L1101 (
	 );
   DFF_X1 L1100 (
	 );
   DFF_X1 L1099 (
	 );
   DFF_X1 L1098 (
	 );
   DFF_X1 L1097 (
	 );
   DFF_X1 L1096 (
	 );
   DFF_X1 L1095 (
	 );
   DFF_X1 L1094 (
	 );
   DFF_X1 L1093 (
	 );
   DFF_X1 L1092 (
	 );
   DFF_X1 L1091 (
	 );
   DFF_X1 L1090 (
	 );
   DFF_X1 L1089 (
	 );
   DFF_X1 L1088 (
	 );
   DFF_X1 L1087 (
	 );
   DFF_X1 L1086 (
	 );
   DFF_X1 L1085 (
	 );
   DFF_X1 L1084 (
	 );
   DFF_X1 L1083 (
	 );
   DFF_X1 L1082 (
	 );
   DFF_X1 L1081 (
	 );
   DFF_X1 L1080 (
	 );
   DFF_X1 L1079 (
	 );
   DFF_X1 L1078 (
	 );
   DFF_X1 L1077 (
	 );
   DFF_X1 L1076 (
	 );
   DFF_X1 L1075 (
	 );
   DFF_X1 L1074 (
	 );
   DFF_X1 L1073 (
	 );
   DFF_X1 L1072 (
	 );
   DFF_X1 L1071 (
	 );
   DFF_X1 L1070 (
	 );
   DFF_X1 L1069 (
	 );
   DFF_X1 L1068 (
	 );
   DFF_X1 L1067 (
	 );
   DFF_X1 L1066 (
	 );
   DFF_X1 L1065 (
	 );
   DFF_X1 L1064 (
	 );
   DFF_X1 L1063 (
	 );
   DFF_X1 L1062 (
	 );
   DFF_X1 L1061 (
	 );
   DFF_X1 L1060 (
	 );
   DFF_X1 L1059 (
	 );
   DFF_X1 L1058 (
	 );
   DFF_X1 L1057 (
	 );
   DFF_X1 L1056 (
	 );
   DFF_X1 L1055 (
	 );
   DFF_X1 L1054 (
	 );
   DFF_X1 L1053 (
	 );
   DFF_X1 L1052 (
	 );
   DFF_X1 L1051 (
	 );
   DFF_X1 L1050 (
	 );
   DFF_X1 L1049 (
	 );
   DFF_X1 L1048 (
	 );
   DFF_X1 L1047 (
	 );
   DFF_X1 L1046 (
	 );
   DFF_X1 L1045 (
	 );
   DFF_X1 L1044 (
	 );
   DFF_X1 L1043 (
	 );
   DFF_X1 L1042 (
	 );
   DFF_X1 L1041 (
	 );
   DFF_X1 L1040 (
	 );
   DFF_X1 L1039 (
	 );
   DFF_X1 L1038 (
	 );
   DFF_X1 L1037 (
	 );
   DFF_X1 L1036 (
	 );
   DFF_X1 L1035 (
	 );
   DFF_X1 L1034 (
	 );
   DFF_X1 L1033 (
	 );
   DFF_X1 L1032 (
	 );
   DFF_X1 L1031 (
	 );
   DFF_X1 L1030 (
	 );
   DFF_X1 L1029 (
	 );
   DFF_X1 L1028 (
	 );
   DFF_X1 L1027 (
	 );
   DFF_X1 L1026 (
	 );
   DFF_X1 L1025 (
	 );
   DFF_X1 L1024 (
	 );
   DFF_X1 L1023 (
	 );
   DFF_X1 L1022 (
	 );
   DFF_X1 L1021 (
	 );
   DFF_X1 L1020 (
	 );
   DFF_X1 L1019 (
	 );
   DFF_X1 L1018 (
	 );
   DFF_X1 L1017 (
	 );
   DFF_X1 L1016 (
	 );
   DFF_X1 L1015 (
	 );
   DFF_X1 L1014 (
	 );
   DFF_X1 L1013 (
	 );
   DFF_X1 L1012 (
	 );
   DFF_X1 L1011 (
	 );
   DFF_X1 L1010 (
	 );
   DFF_X1 L1009 (
	 );
   DFF_X1 L1008 (
	 );
   DFF_X1 L1007 (
	 );
   DFF_X1 L1006 (
	 );
   DFF_X1 L1005 (
	 );
   DFF_X1 L1004 (
	 );
   DFF_X1 L1003 (
	 );
   DFF_X1 L1002 (
	 );
   DFF_X1 L1001 (
	 );
   DFF_X1 L1000 (
	 );
   DFF_X1 L0999 (
	 );
   DFF_X1 L0998 (
	 );
   DFF_X1 L0997 (
	 );
   DFF_X1 L0996 (
	 );
   DFF_X1 L0995 (
	 );
   DFF_X1 L0994 (
	 );
   DFF_X1 L0993 (
	 );
   DFF_X1 L0992 (
	 );
   DFF_X1 L0991 (
	 );
   DFF_X1 L0990 (
	 );
   DFF_X1 L0989 (
	 );
   DFF_X1 L0988 (
	 );
   DFF_X1 L0987 (
	 );
   DFF_X1 L0986 (
	 );
   DFF_X1 L0985 (
	 );
   DFF_X1 L0984 (
	 );
   DFF_X1 L0983 (
	 );
   DFF_X1 L0982 (
	 );
   DFF_X1 L0981 (
	 );
   DFF_X1 L0980 (
	 );
   DFF_X1 L0979 (
	 );
   DFF_X1 L0978 (
	 );
   DFF_X1 L0977 (
	 );
   DFF_X1 L0976 (
	 );
   DFF_X1 L0975 (
	 );
   DFF_X1 L0974 (
	 );
   DFF_X1 L0973 (
	 );
   DFF_X1 L0972 (
	 );
   DFF_X1 L0971 (
	 );
   DFF_X1 L0970 (
	 );
   DFF_X1 L0969 (
	 );
   DFF_X1 L0968 (
	 );
   DFF_X1 L0967 (
	 );
   DFF_X1 L0966 (
	 );
   DFF_X1 L0965 (
	 );
   DFF_X1 L0964 (
	 );
   DFF_X1 L0963 (
	 );
   DFF_X1 L0962 (
	 );
   DFF_X1 L0961 (
	 );
   DFF_X1 L0960 (
	 );
   DFF_X1 L0959 (
	 );
   DFF_X1 L0958 (
	 );
   DFF_X1 L0957 (
	 );
   DFF_X1 L0956 (
	 );
   DFF_X1 L0955 (
	 );
   DFF_X1 L0954 (
	 );
   DFF_X1 L0953 (
	 );
   DFF_X1 L0952 (
	 );
   DFF_X1 L0951 (
	 );
   DFF_X1 L0950 (
	 );
   DFF_X1 L0949 (
	 );
   DFF_X1 L0948 (
	 );
   DFF_X1 L0947 (
	 );
   DFF_X1 L0946 (
	 );
   DFF_X1 L0945 (
	 );
   DFF_X1 L0944 (
	 );
   DFF_X1 L0943 (
	 );
   DFF_X1 L0942 (
	 );
   DFF_X1 L0941 (
	 );
   DFF_X1 L0940 (
	 );
   DFF_X1 L0939 (
	 );
   DFF_X1 L0938 (
	 );
   DFF_X1 L0937 (
	 );
   DFF_X1 L0936 (
	 );
   DFF_X1 L0935 (
	 );
   DFF_X1 L0934 (
	 );
   DFF_X1 L0933 (
	 );
   DFF_X1 L0932 (
	 );
   DFF_X1 L0931 (
	 );
   DFF_X1 L0930 (
	 );
   DFF_X1 L0929 (
	 );
   DFF_X1 L0928 (
	 );
   DFF_X1 L0927 (
	 );
   DFF_X1 L0926 (
	 );
   DFF_X1 L0925 (
	 );
   DFF_X1 L0924 (
	 );
   DFF_X1 L0923 (
	 );
   DFF_X1 L0922 (
	 );
   DFF_X1 L0921 (
	 );
   DFF_X1 L0920 (
	 );
   DFF_X1 L0919 (
	 );
   DFF_X1 L0918 (
	 );
   DFF_X1 L0917 (
	 );
   DFF_X1 L0916 (
	 );
   DFF_X1 L0915 (
	 );
   DFF_X1 L0914 (
	 );
   DFF_X1 L0913 (
	 );
   DFF_X1 L0912 (
	 );
   DFF_X1 L0911 (
	 );
   DFF_X1 L0910 (
	 );
   DFF_X1 L0909 (
	 );
   DFF_X1 L0908 (
	 );
   DFF_X1 L0907 (
	 );
   DFF_X1 L0906 (
	 );
   DFF_X1 L0905 (
	 );
   DFF_X1 L0904 (
	 );
   DFF_X1 L0903 (
	 );
   DFF_X1 L0902 (
	 );
   DFF_X1 L0901 (
	 );
   DFF_X1 L0900 (
	 );
   DFF_X1 L0899 (
	 );
   DFF_X1 L0898 (
	 );
   DFF_X1 L0897 (
	 );
   DFF_X1 L0896 (
	 );
   DFF_X1 L0895 (
	 );
   DFF_X1 L0894 (
	 );
   DFF_X1 L0893 (
	 );
   DFF_X1 L0892 (
	 );
   DFF_X1 L0891 (
	 );
   DFF_X1 L0890 (
	 );
   DFF_X1 L0889 (
	 );
   DFF_X1 L0888 (
	 );
   DFF_X1 L0887 (
	 );
   DFF_X1 L0886 (
	 );
   DFF_X1 L0885 (
	 );
   DFF_X1 L0884 (
	 );
   DFF_X1 L0883 (
	 );
   DFF_X1 L0882 (
	 );
   DFF_X1 L0881 (
	 );
   DFF_X1 L0880 (
	 );
   DFF_X1 L0879 (
	 );
   DFF_X1 L0878 (
	 );
   DFF_X1 L0877 (
	 );
   DFF_X1 L0876 (
	 );
   DFF_X1 L0875 (
	 );
   DFF_X1 L0874 (
	 );
   DFF_X1 L0873 (
	 );
   DFF_X1 L0872 (
	 );
   DFF_X1 L0871 (
	 );
   DFF_X1 L0870 (
	 );
   DFF_X1 L0869 (
	 );
   DFF_X1 L0868 (
	 );
   DFF_X1 L0867 (
	 );
   DFF_X1 L0866 (
	 );
   DFF_X1 L0865 (
	 );
   DFF_X1 L0864 (
	 );
   DFF_X1 L0863 (
	 );
   DFF_X1 L0862 (
	 );
   DFF_X1 L0861 (
	 );
   DFF_X1 L0860 (
	 );
   DFF_X1 L0859 (
	 );
   DFF_X1 L0858 (
	 );
   DFF_X1 L0857 (
	 );
   DFF_X1 L0856 (
	 );
   DFF_X1 L0855 (
	 );
   DFF_X1 L0854 (
	 );
   DFF_X1 L0853 (
	 );
   DFF_X1 L0852 (
	 );
   DFF_X1 L0851 (
	 );
   DFF_X1 L0850 (
	 );
   DFF_X1 L0849 (
	 );
   DFF_X1 L0848 (
	 );
   DFF_X1 L0847 (
	 );
   DFF_X1 L0846 (
	 );
   DFF_X1 L0845 (
	 );
   DFF_X1 L0844 (
	 );
   DFF_X1 L0843 (
	 );
   DFF_X1 L0842 (
	 );
   DFF_X1 L0841 (
	 );
   DFF_X1 L0840 (
	 );
   DFF_X1 L0839 (
	 );
   DFF_X1 L0838 (
	 );
   DFF_X1 L0837 (
	 );
   DFF_X1 L0836 (
	 );
   DFF_X1 L0835 (
	 );
   DFF_X1 L0834 (
	 );
   DFF_X1 L0833 (
	 );
   DFF_X1 L0832 (
	 );
   DFF_X1 L0831 (
	 );
   DFF_X1 L0830 (
	 );
   DFF_X1 L0829 (
	 );
   DFF_X1 L0828 (
	 );
   DFF_X1 L0827 (
	 );
   DFF_X1 L0826 (
	 );
   DFF_X1 L0825 (
	 );
   DFF_X1 L0824 (
	 );
   DFF_X1 L0823 (
	 );
   DFF_X1 L0822 (
	 );
   DFF_X1 L0821 (
	 );
   DFF_X1 L0820 (
	 );
   DFF_X1 L0819 (
	 );
   DFF_X1 L0818 (
	 );
   DFF_X1 L0817 (
	 );
   DFF_X1 L0816 (
	 );
   DFF_X1 L0815 (
	 );
   DFF_X1 L0814 (
	 );
   DFF_X1 L0813 (
	 );
   DFF_X1 L0812 (
	 );
   DFF_X1 L0811 (
	 );
   DFF_X1 L0810 (
	 );
   DFF_X1 L0809 (
	 );
   DFF_X1 L0808 (
	 );
   DFF_X1 L0807 (
	 );
   DFF_X1 L0806 (
	 );
   DFF_X1 L0805 (
	 );
   DFF_X1 L0804 (
	 );
   DFF_X1 L0803 (
	 );
   DFF_X1 L0802 (
	 );
   DFF_X1 L0801 (
	 );
   DFF_X1 L0800 (
	 );
   DFF_X1 L0799 (
	 );
   DFF_X1 L0798 (
	 );
   DFF_X1 L0797 (
	 );
   DFF_X1 L0796 (
	 );
   DFF_X1 L0795 (
	 );
   DFF_X1 L0794 (
	 );
   DFF_X1 L0793 (
	 );
   DFF_X1 L0792 (
	 );
   DFF_X1 L0791 (
	 );
   DFF_X1 L0790 (
	 );
   DFF_X1 L0789 (
	 );
   DFF_X1 L0788 (
	 );
   DFF_X1 L0787 (
	 );
   DFF_X1 L0786 (
	 );
   DFF_X1 L0785 (
	 );
   DFF_X1 L0784 (
	 );
   DFF_X1 L0783 (
	 );
   DFF_X1 L0782 (
	 );
   DFF_X1 L0781 (
	 );
   DFF_X1 L0780 (
	 );
   DFF_X1 L0779 (
	 );
   DFF_X1 L0778 (
	 );
   DFF_X1 L0777 (
	 );
   DFF_X1 L0776 (
	 );
   DFF_X1 L0775 (
	 );
   DFF_X1 L0774 (
	 );
   DFF_X1 L0773 (
	 );
   DFF_X1 L0772 (
	 );
   DFF_X1 L0771 (
	 );
   DFF_X1 L0770 (
	 );
   DFF_X1 L0769 (
	 );
   DFF_X1 L0768 (
	 );
   DFF_X1 L0767 (
	 );
   DFF_X1 L0766 (
	 );
   DFF_X1 L0765 (
	 );
   DFF_X1 L0764 (
	 );
   DFF_X1 L0763 (
	 );
   DFF_X1 L0762 (
	 );
   DFF_X1 L0761 (
	 );
   DFF_X1 L0760 (
	 );
   DFF_X1 L0759 (
	 );
   DFF_X1 L0758 (
	 );
   DFF_X1 L0757 (
	 );
   DFF_X1 L0756 (
	 );
   DFF_X1 L0755 (
	 );
   DFF_X1 L0754 (
	 );
   DFF_X1 L0753 (
	 );
   DFF_X1 L0752 (
	 );
   DFF_X1 L0751 (
	 );
   DFF_X1 L0750 (
	 );
   DFF_X1 L0749 (
	 );
   DFF_X1 L0748 (
	 );
   DFF_X1 L0747 (
	 );
   DFF_X1 L0746 (
	 );
   DFF_X1 L0745 (
	 );
   DFF_X1 L0744 (
	 );
   DFF_X1 L0743 (
	 );
   DFF_X1 L0742 (
	 );
   DFF_X1 L0741 (
	 );
   DFF_X1 L0740 (
	 );
   DFF_X1 L0739 (
	 );
   DFF_X1 L0738 (
	 );
   DFF_X1 L0737 (
	 );
   DFF_X1 L0736 (
	 );
   DFF_X1 L0735 (
	 );
   DFF_X1 L0734 (
	 );
   DFF_X1 L0733 (
	 );
   DFF_X1 L0732 (
	 );
   DFF_X1 L0731 (
	 );
   DFF_X1 L0730 (
	 );
   DFF_X1 L0729 (
	 );
   DFF_X1 L0728 (
	 );
   DFF_X1 L0727 (
	 );
   DFF_X1 L0726 (
	 );
   DFF_X1 L0725 (
	 );
   DFF_X1 L0724 (
	 );
   DFF_X1 L0723 (
	 );
   DFF_X1 L0722 (
	 );
   DFF_X1 L0721 (
	 );
   DFF_X1 L0720 (
	 );
   DFF_X1 L0719 (
	 );
   DFF_X1 L0718 (
	 );
   DFF_X1 L0717 (
	 );
   DFF_X1 L0716 (
	 );
   DFF_X1 L0715 (
	 );
   DFF_X1 L0714 (
	 );
   DFF_X1 L0713 (
	 );
   DFF_X1 L0712 (
	 );
   DFF_X1 L0711 (
	 );
   DFF_X1 L0710 (
	 );
   DFF_X1 L0709 (
	 );
   DFF_X1 L0708 (
	 );
   DFF_X1 L0707 (
	 );
   DFF_X1 L0706 (
	 );
   DFF_X1 L0705 (
	 );
   DFF_X1 L0704 (
	 );
   DFF_X1 L0703 (
	 );
   DFF_X1 L0702 (
	 );
   DFF_X1 L0701 (
	 );
   DFF_X1 L0700 (
	 );
   DFF_X1 L0699 (
	 );
   DFF_X1 L0698 (
	 );
   DFF_X1 L0697 (
	 );
   DFF_X1 L0696 (
	 );
   DFF_X1 L0695 (
	 );
   DFF_X1 L0694 (
	 );
   DFF_X1 L0693 (
	 );
   DFF_X1 L0692 (
	 );
   DFF_X1 L0691 (
	 );
   DFF_X1 L0690 (
	 );
   DFF_X1 L0689 (
	 );
   DFF_X1 L0688 (
	 );
   DFF_X1 L0687 (
	 );
   DFF_X1 L0686 (
	 );
   DFF_X1 L0685 (
	 );
   DFF_X1 L0684 (
	 );
   DFF_X1 L0683 (
	 );
   DFF_X1 L0682 (
	 );
   DFF_X1 L0681 (
	 );
   DFF_X1 L0680 (
	 );
   DFF_X1 L0679 (
	 );
   DFF_X1 L0678 (
	 );
   DFF_X1 L0677 (
	 );
   DFF_X1 L0676 (
	 );
   DFF_X1 L0675 (
	 );
   DFF_X1 L0674 (
	 );
   DFF_X1 L0673 (
	 );
   DFF_X1 L0672 (
	 );
   DFF_X1 L0671 (
	 );
   DFF_X1 L0670 (
	 );
   DFF_X1 L0669 (
	 );
   DFF_X1 L0668 (
	 );
   DFF_X1 L0667 (
	 );
   DFF_X1 L0666 (
	 );
   DFF_X1 L0665 (
	 );
   DFF_X1 L0664 (
	 );
   DFF_X1 L0663 (
	 );
   DFF_X1 L0662 (
	 );
   DFF_X1 L0661 (
	 );
   DFF_X1 L0660 (
	 );
   DFF_X1 L0659 (
	 );
   DFF_X1 L0658 (
	 );
   DFF_X1 L0657 (
	 );
   DFF_X1 L0656 (
	 );
   DFF_X1 L0655 (
	 );
   DFF_X1 L0654 (
	 );
   DFF_X1 L0653 (
	 );
   DFF_X1 L0652 (
	 );
   DFF_X1 L0651 (
	 );
   DFF_X1 L0650 (
	 );
   DFF_X1 L0649 (
	 );
   DFF_X1 L0648 (
	 );
   DFF_X1 L0647 (
	 );
   DFF_X1 L0646 (
	 );
   DFF_X1 L0645 (
	 );
   DFF_X1 L0644 (
	 );
   DFF_X1 L0643 (
	 );
   DFF_X1 L0642 (
	 );
   DFF_X1 L0641 (
	 );
   DFF_X1 L0640 (
	 );
   DFF_X1 L0639 (
	 );
   DFF_X1 L0638 (
	 );
   DFF_X1 L0637 (
	 );
   DFF_X1 L0636 (
	 );
   DFF_X1 L0635 (
	 );
   DFF_X1 L0634 (
	 );
   DFF_X1 L0633 (
	 );
   DFF_X1 L0632 (
	 );
   DFF_X1 L0631 (
	 );
   DFF_X1 L0630 (
	 );
   DFF_X1 L0629 (
	 );
   DFF_X1 L0628 (
	 );
   DFF_X1 L0627 (
	 );
   DFF_X1 L0626 (
	 );
   DFF_X1 L0625 (
	 );
   DFF_X1 L0624 (
	 );
   DFF_X1 L0623 (
	 );
   DFF_X1 L0622 (
	 );
   DFF_X1 L0621 (
	 );
   DFF_X1 L0620 (
	 );
   DFF_X1 L0619 (
	 );
   DFF_X1 L0618 (
	 );
   DFF_X1 L0617 (
	 );
   DFF_X1 L0616 (
	 );
   DFF_X1 L0615 (
	 );
   DFF_X1 L0614 (
	 );
   DFF_X1 L0613 (
	 );
   DFF_X1 L0612 (
	 );
   DFF_X1 L0611 (
	 );
   DFF_X1 L0610 (
	 );
   DFF_X1 L0609 (
	 );
   DFF_X1 L0608 (
	 );
   DFF_X1 L0607 (
	 );
   DFF_X1 L0606 (
	 );
   DFF_X1 L0605 (
	 );
   DFF_X1 L0604 (
	 );
   DFF_X1 L0603 (
	 );
   DFF_X1 L0602 (
	 );
   DFF_X1 L0601 (
	 );
   DFF_X1 L0600 (
	 );
   DFF_X1 L0599 (
	 );
   DFF_X1 L0598 (
	 );
   DFF_X1 L0597 (
	 );
   DFF_X1 L0596 (
	 );
   DFF_X1 L0595 (
	 );
   DFF_X1 L0594 (
	 );
   DFF_X1 L0593 (
	 );
   DFF_X1 L0592 (
	 );
   DFF_X1 L0591 (
	 );
   DFF_X1 L0590 (
	 );
   DFF_X1 L0589 (
	 );
   DFF_X1 L0588 (
	 );
   DFF_X1 L0587 (
	 );
   DFF_X1 L0586 (
	 );
   DFF_X1 L0585 (
	 );
   DFF_X1 L0584 (
	 );
   DFF_X1 L0583 (
	 );
   DFF_X1 L0582 (
	 );
   DFF_X1 L0581 (
	 );
   DFF_X1 L0580 (
	 );
   DFF_X1 L0579 (
	 );
   DFF_X1 L0578 (
	 );
   DFF_X1 L0577 (
	 );
   DFF_X1 L0576 (
	 );
   DFF_X1 L0575 (
	 );
   DFF_X1 L0574 (
	 );
   DFF_X1 L0573 (
	 );
   DFF_X1 L0572 (
	 );
   DFF_X1 L0571 (
	 );
   DFF_X1 L0570 (
	 );
   DFF_X1 L0569 (
	 );
   DFF_X1 L0568 (
	 );
   DFF_X1 L0567 (
	 );
   DFF_X1 L0566 (
	 );
   DFF_X1 L0565 (
	 );
   DFF_X1 L0564 (
	 );
   DFF_X1 L0563 (
	 );
   DFF_X1 L0562 (
	 );
   DFF_X1 L0561 (
	 );
   DFF_X1 L0560 (
	 );
   DFF_X1 L0559 (
	 );
   DFF_X1 L0558 (
	 );
   DFF_X1 L0557 (
	 );
   DFF_X1 L0556 (
	 );
   DFF_X1 L0555 (
	 );
   DFF_X1 L0554 (
	 );
   DFF_X1 L0553 (
	 );
   DFF_X1 L0552 (
	 );
   DFF_X1 L0551 (
	 );
   DFF_X1 L0550 (
	 );
   DFF_X1 L0549 (
	 );
   DFF_X1 L0548 (
	 );
   DFF_X1 L0547 (
	 );
   DFF_X1 L0546 (
	 );
   DFF_X1 L0545 (
	 );
   DFF_X1 L0544 (
	 );
   DFF_X1 L0543 (
	 );
   DFF_X1 L0542 (
	 );
   DFF_X1 L0541 (
	 );
   DFF_X1 L0540 (
	 );
   DFF_X1 L0539 (
	 );
   DFF_X1 L0538 (
	 );
   DFF_X1 L0537 (
	 );
   DFF_X1 L0536 (
	 );
   DFF_X1 L0535 (
	 );
   DFF_X1 L0534 (
	 );
   DFF_X1 L0533 (
	 );
   DFF_X1 L0532 (
	 );
   DFF_X1 L0531 (
	 );
   DFF_X1 L0530 (
	 );
   DFF_X1 L0529 (
	 );
   DFF_X1 L0528 (
	 );
   DFF_X1 L0527 (
	 );
   DFF_X1 L0526 (
	 );
   DFF_X1 L0525 (
	 );
   DFF_X1 L0524 (
	 );
   DFF_X1 L0523 (
	 );
   DFF_X1 L0522 (
	 );
   DFF_X1 L0521 (
	 );
   DFF_X1 L0520 (
	 );
   DFF_X1 L0519 (
	 );
   DFF_X1 L0518 (
	 );
   DFF_X1 L0517 (
	 );
   DFF_X1 L0516 (
	 );
   DFF_X1 L0515 (
	 );
   DFF_X1 L0514 (
	 );
   DFF_X1 L0513 (
	 );
   DFF_X1 L0512 (
	 );
   DFF_X1 L0511 (
	 );
   DFF_X1 L0510 (
	 );
   DFF_X1 L0509 (
	 );
   DFF_X1 L0508 (
	 );
   DFF_X1 L0507 (
	 );
   DFF_X1 L0506 (
	 );
   DFF_X1 L0505 (
	 );
   DFF_X1 L0504 (
	 );
   DFF_X1 L0503 (
	 );
   DFF_X1 L0502 (
	 );
   DFF_X1 L0501 (
	 );
   DFF_X1 L0500 (
	 );
   DFF_X1 L0499 (
	 );
   DFF_X1 L0498 (
	 );
   DFF_X1 L0497 (
	 );
   DFF_X1 L0496 (
	 );
   DFF_X1 L0495 (
	 );
   DFF_X1 L0494 (
	 );
   DFF_X1 L0493 (
	 );
   DFF_X1 L0492 (
	 );
   DFF_X1 L0491 (
	 );
   DFF_X1 L0490 (
	 );
   DFF_X1 L0489 (
	 );
   DFF_X1 L0488 (
	 );
   DFF_X1 L0487 (
	 );
   DFF_X1 L0486 (
	 );
   DFF_X1 L0485 (
	 );
   DFF_X1 L0484 (
	 );
   DFF_X1 L0483 (
	 );
   DFF_X1 L0482 (
	 );
   DFF_X1 L0481 (
	 );
   DFF_X1 L0480 (
	 );
   DFF_X1 L0479 (
	 );
   DFF_X1 L0478 (
	 );
   DFF_X1 L0477 (
	 );
   DFF_X1 L0476 (
	 );
   DFF_X1 L0475 (
	 );
   DFF_X1 L0474 (
	 );
   DFF_X1 L0473 (
	 );
   DFF_X1 L0472 (
	 );
   DFF_X1 L0471 (
	 );
   DFF_X1 L0470 (
	 );
   DFF_X1 L0469 (
	 );
   DFF_X1 L0468 (
	 );
   DFF_X1 L0467 (
	 );
   DFF_X1 L0466 (
	 );
   DFF_X1 L0465 (
	 );
   DFF_X1 L0464 (
	 );
   DFF_X1 L0463 (
	 );
   DFF_X1 L0462 (
	 );
   DFF_X1 L0461 (
	 );
   DFF_X1 L0460 (
	 );
   DFF_X1 L0459 (
	 );
   DFF_X1 L0458 (
	 );
   DFF_X1 L0457 (
	 );
   DFF_X1 L0456 (
	 );
   DFF_X1 L0455 (
	 );
   DFF_X1 L0454 (
	 );
   DFF_X1 L0453 (
	 );
   DFF_X1 L0452 (
	 );
   DFF_X1 L0451 (
	 );
   DFF_X1 L0450 (
	 );
   DFF_X1 L0449 (
	 );
   DFF_X1 L0448 (
	 );
   DFF_X1 L0447 (
	 );
   DFF_X1 L0446 (
	 );
   DFF_X1 L0445 (
	 );
   DFF_X1 L0444 (
	 );
   DFF_X1 L0443 (
	 );
   DFF_X1 L0442 (
	 );
   DFF_X1 L0441 (
	 );
   DFF_X1 L0440 (
	 );
   DFF_X1 L0439 (
	 );
   DFF_X1 L0438 (
	 );
   DFF_X1 L0437 (
	 );
   DFF_X1 L0436 (
	 );
   DFF_X1 L0435 (
	 );
   DFF_X1 L0434 (
	 );
   DFF_X1 L0433 (
	 );
   DFF_X1 L0432 (
	 );
   DFF_X1 L0431 (
	 );
   DFF_X1 L0430 (
	 );
   DFF_X1 L0429 (
	 );
   DFF_X1 L0428 (
	 );
   DFF_X1 L0427 (
	 );
   DFF_X1 L0426 (
	 );
   DFF_X1 L0425 (
	 );
   DFF_X1 L0424 (
	 );
   DFF_X1 L0423 (
	 );
   DFF_X1 L0422 (
	 );
   DFF_X1 L0421 (
	 );
   DFF_X1 L0420 (
	 );
   DFF_X1 L0419 (
	 );
   DFF_X1 L0418 (
	 );
   DFF_X1 L0417 (
	 );
   DFF_X1 L0416 (
	 );
   DFF_X1 L0415 (
	 );
   DFF_X1 L0414 (
	 );
   DFF_X1 L0413 (
	 );
   DFF_X1 L0412 (
	 );
   DFF_X1 L0411 (
	 );
   DFF_X1 L0410 (
	 );
   DFF_X1 L0409 (
	 );
   DFF_X1 L0408 (
	 );
   DFF_X1 L0407 (
	 );
   DFF_X1 L0406 (
	 );
   DFF_X1 L0405 (
	 );
   DFF_X1 L0404 (
	 );
   DFF_X1 L0403 (
	 );
   DFF_X1 L0402 (
	 );
   DFF_X1 L0401 (
	 );
   DFF_X1 L0400 (
	 );
   DFF_X1 L0399 (
	 );
   DFF_X1 L0398 (
	 );
   DFF_X1 L0397 (
	 );
   DFF_X1 L0396 (
	 );
   DFF_X1 L0395 (
	 );
   DFF_X1 L0394 (
	 );
   DFF_X1 L0393 (
	 );
   DFF_X1 L0392 (
	 );
   DFF_X1 L0391 (
	 );
   DFF_X1 L0390 (
	 );
   DFF_X1 L0389 (
	 );
   DFF_X1 L0388 (
	 );
   DFF_X1 L0387 (
	 );
   DFF_X1 L0386 (
	 );
   DFF_X1 L0385 (
	 );
   DFF_X1 L0384 (
	 );
   DFF_X1 L0383 (
	 );
   DFF_X1 L0382 (
	 );
   DFF_X1 L0381 (
	 );
   DFF_X1 L0380 (
	 );
   DFF_X1 L0379 (
	 );
   DFF_X1 L0378 (
	 );
   DFF_X1 L0377 (
	 );
   DFF_X1 L0376 (
	 );
   DFF_X1 L0375 (
	 );
   DFF_X1 L0374 (
	 );
   DFF_X1 L0373 (
	 );
   DFF_X1 L0372 (
	 );
   DFF_X1 L0371 (
	 );
   DFF_X1 L0370 (
	 );
   DFF_X1 L0369 (
	 );
   DFF_X1 L0368 (
	 );
   DFF_X1 L0367 (
	 );
   DFF_X1 L0366 (
	 );
   DFF_X1 L0365 (
	 );
   DFF_X1 L0364 (
	 );
   DFF_X1 L0363 (
	 );
   DFF_X1 L0362 (
	 );
   DFF_X1 L0361 (
	 );
   DFF_X1 L0360 (
	 );
   DFF_X1 L0359 (
	 );
   DFF_X1 L0358 (
	 );
   DFF_X1 L0357 (
	 );
   DFF_X1 L0356 (
	 );
   DFF_X1 L0355 (
	 );
   DFF_X1 L0354 (
	 );
   DFF_X1 L0353 (
	 );
   DFF_X1 L0352 (
	 );
   DFF_X1 L0351 (
	 );
   DFF_X1 L0350 (
	 );
   DFF_X1 L0349 (
	 );
   DFF_X1 L0348 (
	 );
   DFF_X1 L0347 (
	 );
   DFF_X1 L0346 (
	 );
   DFF_X1 L0345 (
	 );
   DFF_X1 L0344 (
	 );
   DFF_X1 L0343 (
	 );
   DFF_X1 L0342 (
	 );
   DFF_X1 L0341 (
	 );
   DFF_X1 L0340 (
	 );
   DFF_X1 L0339 (
	 );
   DFF_X1 L0338 (
	 );
   DFF_X1 L0337 (
	 );
   DFF_X1 L0336 (
	 );
   DFF_X1 L0335 (
	 );
   DFF_X1 L0334 (
	 );
   DFF_X1 L0333 (
	 );
   DFF_X1 L0332 (
	 );
   DFF_X1 L0331 (
	 );
   DFF_X1 L0330 (
	 );
   DFF_X1 L0329 (
	 );
   DFF_X1 L0328 (
	 );
   DFF_X1 L0327 (
	 );
   DFF_X1 L0326 (
	 );
   DFF_X1 L0325 (
	 );
   DFF_X1 L0324 (
	 );
   DFF_X1 L0323 (
	 );
   DFF_X1 L0322 (
	 );
   DFF_X1 L0321 (
	 );
   DFF_X1 L0320 (
	 );
   DFF_X1 L0319 (
	 );
   DFF_X1 L0318 (
	 );
   DFF_X1 L0317 (
	 );
   DFF_X1 L0316 (
	 );
   DFF_X1 L0315 (
	 );
   DFF_X1 L0314 (
	 );
   DFF_X1 L0313 (
	 );
   DFF_X1 L0312 (
	 );
   DFF_X1 L0311 (
	 );
   DFF_X1 L0310 (
	 );
   DFF_X1 L0309 (
	 );
   DFF_X1 L0308 (
	 );
   DFF_X1 L0307 (
	 );
   DFF_X1 L0306 (
	 );
   DFF_X1 L0305 (
	 );
   DFF_X1 L0304 (
	 );
   DFF_X1 L0303 (
	 );
   DFF_X1 L0302 (
	 );
   DFF_X1 L0301 (
	 );
   DFF_X1 L0300 (
	 );
   DFF_X1 L0299 (
	 );
   DFF_X1 L0298 (
	 );
   DFF_X1 L0297 (
	 );
   DFF_X1 L0296 (
	 );
   DFF_X1 L0295 (
	 );
   DFF_X1 L0294 (
	 );
   DFF_X1 L0293 (
	 );
   DFF_X1 L0292 (
	 );
   DFF_X1 L0291 (
	 );
   DFF_X1 L0290 (
	 );
   DFF_X1 L0289 (
	 );
   DFF_X1 L0288 (
	 );
   DFF_X1 L0287 (
	 );
   DFF_X1 L0286 (
	 );
   DFF_X1 L0285 (
	 );
   DFF_X1 L0284 (
	 );
   DFF_X1 L0283 (
	 );
   DFF_X1 L0282 (
	 );
   DFF_X1 L0281 (
	 );
   DFF_X1 L0280 (
	 );
   DFF_X1 L0279 (
	 );
   DFF_X1 L0278 (
	 );
   DFF_X1 L0277 (
	 );
   DFF_X1 L0276 (
	 );
   DFF_X1 L0275 (
	 );
   DFF_X1 L0274 (
	 );
   DFF_X1 L0273 (
	 );
   DFF_X1 L0272 (
	 );
   DFF_X1 L0271 (
	 );
   DFF_X1 L0270 (
	 );
   DFF_X1 L0269 (
	 );
   DFF_X1 L0268 (
	 );
   DFF_X1 L0267 (
	 );
   DFF_X1 L0266 (
	 );
   DFF_X1 L0265 (
	 );
   DFF_X1 L0264 (
	 );
   DFF_X1 L0263 (
	 );
   DFF_X1 L0262 (
	 );
   DFF_X1 L0261 (
	 );
   DFF_X1 L0260 (
	 );
   DFF_X1 L0259 (
	 );
   DFF_X1 L0258 (
	 );
   DFF_X1 L0257 (
	 );
   DFF_X1 L0256 (
	 );
   DFF_X1 L0255 (
	 );
   DFF_X1 L0254 (
	 );
   DFF_X1 L0253 (
	 );
   DFF_X1 L0252 (
	 );
   DFF_X1 L0251 (
	 );
   DFF_X1 L0250 (
	 );
   DFF_X1 L0249 (
	 );
   DFF_X1 L0248 (
	 );
   DFF_X1 L0247 (
	 );
   DFF_X1 L0246 (
	 );
   DFF_X1 L0245 (
	 );
   DFF_X1 L0244 (
	 );
   DFF_X1 L0243 (
	 );
   DFF_X1 L0242 (
	 );
   DFF_X1 L0241 (
	 );
   DFF_X1 L0240 (
	 );
   DFF_X1 L0239 (
	 );
   DFF_X1 L0238 (
	 );
   DFF_X1 L0237 (
	 );
   DFF_X1 L0236 (
	 );
   DFF_X1 L0235 (
	 );
   DFF_X1 L0234 (
	 );
   DFF_X1 L0233 (
	 );
   DFF_X1 L0232 (
	 );
   DFF_X1 L0231 (
	 );
   DFF_X1 L0230 (
	 );
   DFF_X1 L0229 (
	 );
   DFF_X1 L0228 (
	 );
   DFF_X1 L0227 (
	 );
   DFF_X1 L0226 (
	 );
   DFF_X1 L0225 (
	 );
   DFF_X1 L0224 (
	 );
   DFF_X1 L0223 (
	 );
   DFF_X1 L0222 (
	 );
   DFF_X1 L0221 (
	 );
   DFF_X1 L0220 (
	 );
   DFF_X1 L0219 (
	 );
   DFF_X1 L0218 (
	 );
   DFF_X1 L0217 (
	 );
   DFF_X1 L0216 (
	 );
   DFF_X1 L0215 (
	 );
   DFF_X1 L0214 (
	 );
   DFF_X1 L0213 (
	 );
   DFF_X1 L0212 (
	 );
   DFF_X1 L0211 (
	 );
   DFF_X1 L0210 (
	 );
   DFF_X1 L0209 (
	 );
   DFF_X1 L0208 (
	 );
   DFF_X1 L0207 (
	 );
   DFF_X1 L0206 (
	 );
   DFF_X1 L0205 (
	 );
   DFF_X1 L0204 (
	 );
   DFF_X1 L0203 (
	 );
   DFF_X1 L0202 (
	 );
   DFF_X1 L0201 (
	 );
   DFF_X1 L0200 (
	 );
   DFF_X1 L0199 (
	 );
   DFF_X1 L0198 (
	 );
   DFF_X1 L0197 (
	 );
   DFF_X1 L0196 (
	 );
   DFF_X1 L0195 (
	 );
   DFF_X1 L0194 (
	 );
   DFF_X1 L0193 (
	 );
   DFF_X1 L0192 (
	 );
   DFF_X1 L0191 (
	 );
   DFF_X1 L0190 (
	 );
   DFF_X1 L0189 (
	 );
   DFF_X1 L0188 (
	 );
   DFF_X1 L0187 (
	 );
   DFF_X1 L0186 (
	 );
   DFF_X1 L0185 (
	 );
   DFF_X1 L0184 (
	 );
   DFF_X1 L0183 (
	 );
   DFF_X1 L0182 (
	 );
   DFF_X1 L0181 (
	 );
   DFF_X1 L0180 (
	 );
   DFF_X1 L0179 (
	 );
   DFF_X1 L0178 (
	 );
   DFF_X1 L0177 (
	 );
   DFF_X1 L0176 (
	 );
   DFF_X1 L0175 (
	 );
   DFF_X1 L0174 (
	 );
   DFF_X1 L0173 (
	 );
   DFF_X1 L0172 (
	 );
   DFF_X1 L0171 (
	 );
   DFF_X1 L0170 (
	 );
   DFF_X1 L0169 (
	 );
   DFF_X1 L0168 (
	 );
   DFF_X1 L0167 (
	 );
   DFF_X1 L0166 (
	 );
   DFF_X1 L0165 (
	 );
   DFF_X1 L0164 (
	 );
   DFF_X1 L0163 (
	 );
   DFF_X1 L0162 (
	 );
   DFF_X1 L0161 (
	 );
   DFF_X1 L0160 (
	 );
   DFF_X1 L0159 (
	 );
   DFF_X1 L0158 (
	 );
   DFF_X1 L0157 (
	 );
   DFF_X1 L0156 (
	 );
   DFF_X1 L0155 (
	 );
   DFF_X1 L0154 (
	 );
   DFF_X1 L0153 (
	 );
   DFF_X1 L0152 (
	 );
   DFF_X1 L0151 (
	 );
   DFF_X1 L0150 (
	 );
   DFF_X1 L0149 (
	 );
   DFF_X1 L0148 (
	 );
   DFF_X1 L0147 (
	 );
   DFF_X1 L0146 (
	 );
   DFF_X1 L0145 (
	 );
   DFF_X1 L0144 (
	 );
   DFF_X1 L0143 (
	 );
   DFF_X1 L0142 (
	 );
   DFF_X1 L0141 (
	 );
   DFF_X1 L0140 (
	 );
   DFF_X1 L0139 (
	 );
   DFF_X1 L0138 (
	 );
   DFF_X1 L0137 (
	 );
   DFF_X1 L0136 (
	 );
   DFF_X1 L0135 (
	 );
   DFF_X1 L0134 (
	 );
   DFF_X1 L0133 (
	 );
   DFF_X1 L0132 (
	 );
   DFF_X1 L0131 (
	 );
   DFF_X1 L0130 (
	 );
   DFF_X1 L0129 (
	 );
   DFF_X1 L0128 (
	 );
   DFF_X1 L0127 (
	 );
   DFF_X1 L0126 (
	 );
   DFF_X1 L0125 (
	 );
   DFF_X1 L0124 (
	 );
   DFF_X1 L0123 (
	 );
   DFF_X1 L0122 (
	 );
   DFF_X1 L0121 (
	 );
   DFF_X1 L0120 (
	 );
   DFF_X1 L0119 (
	 );
   DFF_X1 L0118 (
	 );
   DFF_X1 L0117 (
	 );
   DFF_X1 L0116 (
	 );
   DFF_X1 L0115 (
	 );
   DFF_X1 L0114 (
	 );
   DFF_X1 L0113 (
	 );
   DFF_X1 L0112 (
	 );
   DFF_X1 L0111 (
	 );
   DFF_X1 L0110 (
	 );
   DFF_X1 L0109 (
	 );
   DFF_X1 L0108 (
	 );
   DFF_X1 L0107 (
	 );
   DFF_X1 L0106 (
	 );
   DFF_X1 L0105 (
	 );
   DFF_X1 L0104 (
	 );
   DFF_X1 L0103 (
	 );
   DFF_X1 L0102 (
	 );
   DFF_X1 L0101 (
	 );
   DFF_X1 L0100 (
	 );
   DFF_X1 L0099 (
	 );
   DFF_X1 L0098 (
	 );
   DFF_X1 L0097 (
	 );
   DFF_X1 L0096 (
	 );
   DFF_X1 L0095 (
	 );
   DFF_X1 L0094 (
	 );
   DFF_X1 L0093 (
	 );
   DFF_X1 L0092 (
	 );
   DFF_X1 L0091 (
	 );
   DFF_X1 L0090 (
	 );
   DFF_X1 L0089 (
	 );
   DFF_X1 L0088 (
	 );
   DFF_X1 L0087 (
	 );
   DFF_X1 L0086 (
	 );
   DFF_X1 L0085 (
	 );
   DFF_X1 L0084 (
	 );
   DFF_X1 L0083 (
	 );
   DFF_X1 L0082 (
	 );
   DFF_X1 L0081 (
	 );
   DFF_X1 L0080 (
	 );
   DFF_X1 L0079 (
	 );
   DFF_X1 L0078 (
	 );
   DFF_X1 L0077 (
	 );
   DFF_X1 L0076 (
	 );
   DFF_X1 L0075 (
	 );
   DFF_X1 L0074 (
	 );
   DFF_X1 L0073 (
	 );
   DFF_X1 L0072 (
	 );
   DFF_X1 L0071 (
	 );
   DFF_X1 L0070 (
	 );
   DFF_X1 L0069 (
	 );
   DFF_X1 L0068 (
	 );
   DFF_X1 L0067 (
	 );
   DFF_X1 L0066 (
	 );
   DFF_X1 L0065 (
	 );
   DFF_X1 L0064 (
	 );
   DFF_X1 L0063 (
	 );
   DFF_X1 L0062 (
	 );
   DFF_X1 L0061 (
	 );
   DFF_X1 L0060 (
	 );
   DFF_X1 L0059 (
	 );
   DFF_X1 L0058 (
	 );
   DFF_X1 L0057 (
	 );
   DFF_X1 L0056 (
	 );
   DFF_X1 L0055 (
	 );
   DFF_X1 L0054 (
	 );
   DFF_X1 L0053 (
	 );
   DFF_X1 L0052 (
	 );
   DFF_X1 L0051 (
	 );
   DFF_X1 L0050 (
	 );
   DFF_X1 L0049 (
	 );
   DFF_X1 L0048 (
	 );
   DFF_X1 L0047 (
	 );
   DFF_X1 L0046 (
	 );
   DFF_X1 L0045 (
	 );
   DFF_X1 L0044 (
	 );
   DFF_X1 L0043 (
	 );
   DFF_X1 L0042 (
	 );
   DFF_X1 L0041 (
	 );
   DFF_X1 L0040 (
	 );
   DFF_X1 L0039 (
	 );
   DFF_X1 L0038 (
	 );
   DFF_X1 L0037 (
	 );
   DFF_X1 L0036 (
	 );
   DFF_X1 L0035 (
	 );
   DFF_X1 L0034 (
	 );
   DFF_X1 L0033 (
	 );
   DFF_X1 L0032 (
	 );
   DFF_X1 L0031 (
	 );
   DFF_X1 L0030 (
	 );
   DFF_X1 L0029 (
	 );
   DFF_X1 L0028 (
	 );
   DFF_X1 L0027 (
	 );
   DFF_X1 L0026 (
	 );
   DFF_X1 L0025 (
	 );
   DFF_X1 L0024 (
	 );
   DFF_X1 L0023 (
	 );
   DFF_X1 L0022 (
	 );
   DFF_X1 L0021 (
	 );
   DFF_X1 L0020 (
	 );
   DFF_X1 L0019 (
	 );
   DFF_X1 L0018 (
	 );
   DFF_X1 L0017 (
	 );
   DFF_X1 L0016 (
	 );
   DFF_X1 L0015 (
	 );
   DFF_X1 L0014 (
	 );
   DFF_X1 L0013 (
	 );
   DFF_X1 L0012 (
	 );
   DFF_X1 L0011 (
	 );
   DFF_X1 L0010 (
	 );
   DFF_X1 L0009 (
	 );
   DFF_X1 L0008 (
	 );
   DFF_X1 L0007 (
	 );
   DFF_X1 L0006 (
	 );
   DFF_X1 L0005 (
	 );
   DFF_X1 L0004 (
	 );
   DFF_X1 L0003 (
	 );
   DFF_X1 L0002 (
	 );
   DFF_X1 L0001 (
	 );
   CLKBUF_X1 G5608 (
	 );
   CLKBUF_X1 G5607 (
	 );
   OAI21_X1 G5606 (
	 );
   NAND2_X1 G5605 (
	 );
   NOR2_X1 G5604 (
	 );
   CLKBUF_X1 G5603 (
	 );
   NAND3_X1 G5602 (
	 );
   AOI22_X1 G5601 (
	 );
   AND3_X1 G5600 (
	 );
   NAND2_X1 G5599 (
	 );
   NAND2_X1 G5598 (
	 );
   NAND2_X1 G5597 (
	 );
   AND3_X1 G5596 (
	 );
   NAND4_X1 G5595 (
	 );
   NAND4_X1 G5594 (
	 );
   NAND4_X1 G5593 (
	 );
   CLKBUF_X1 G5592 (
	 );
   OAI21_X1 G5591 (
	 );
   NAND2_X1 G5590 (
	 );
   CLKBUF_X1 G5589 (
	 );
   CLKBUF_X1 G5588 (
	 );
   NAND2_X1 G5587 (
	 );
   AOI22_X1 G5586 (
	 );
   AOI22_X1 G5585 (
	 );
   CLKBUF_X1 G5584 (
	 );
   CLKBUF_X1 G5583 (
	 );
   CLKBUF_X1 G5582 (
	 );
   OAI21_X1 G5581 (
	 );
   NAND2_X1 G5580 (
	 );
   OAI21_X1 G5579 (
	 );
   INV_X1 G5578 (
	 );
   NAND2_X1 G5577 (
	 );
   NAND3_X1 G5576 (
	 );
   AOI22_X1 G5575 (
	 );
   AND3_X1 G5574 (
	 );
   NAND2_X1 G5573 (
	 );
   NAND2_X1 G5572 (
	 );
   NAND2_X1 G5571 (
	 );
   AND3_X1 G5570 (
	 );
   NAND4_X1 G5569 (
	 );
   NAND4_X1 G5568 (
	 );
   NAND4_X1 G5567 (
	 );
   NAND4_X1 G5566 (
	 );
   AOI22_X1 G5565 (
	 );
   NAND2_X1 G5564 (
	 );
   NAND2_X1 G5563 (
	 );
   NAND2_X1 G5562 (
	 );
   OAI211_X1 G5561 (
	 );
   INV_X1 G5560 (
	 );
   NAND2_X1 G5559 (
	 );
   OAI21_X1 G5558 (
	 );
   OAI21_X1 G5557 (
	 );
   INV_X1 G5556 (
	 );
   NAND2_X1 G5555 (
	 );
   CLKBUF_X1 G5554 (
	 );
   NAND3_X1 G5553 (
	 );
   OR2_X1 G5552 (
	 );
   NOR3_X1 G5551 (
	 );
   NAND3_X1 G5550 (
	 );
   NAND4_X1 G5549 (
	 );
   NAND3_X1 G5548 (
	 );
   NAND3_X1 G5547 (
	 );
   OAI22_X1 G5546 (
	 );
   INV_X1 G5545 (
	 );
   AND4_X1 G5544 (
	 );
   NOR2_X1 G5543 (
	 );
   NOR2_X1 G5542 (
	 );
   NOR2_X1 G5541 (
	 );
   INV_X1 G5540 (
	 );
   NOR2_X1 G5539 (
	 );
   NAND2_X1 G5538 (
	 );
   AND2_X1 G5537 (
	 );
   OAI21_X1 G5536 (
	 );
   NAND2_X1 G5535 (
	 );
   CLKBUF_X1 G5534 (
	 );
   AND2_X1 G5533 (
	 );
   MUX2_X1 G5532 (
	 );
   MUX2_X1 G5531 (
	 );
   CLKBUF_X1 G5530 (
	 );
   CLKBUF_X1 G5529 (
	 );
   MUX2_X1 G5528 (
	 );
   CLKBUF_X1 G5527 (
	 );
   CLKBUF_X1 G5526 (
	 );
   CLKBUF_X1 G5525 (
	 );
   CLKBUF_X1 G5524 (
	 );
   MUX2_X1 G5523 (
	 );
   CLKBUF_X1 G5522 (
	 );
   CLKBUF_X1 G5521 (
	 );
   CLKBUF_X1 G5520 (
	 );
   NOR3_X1 G5519 (
	 );
   NOR2_X1 G5518 (
	 );
   CLKBUF_X1 G5517 (
	 );
   NAND3_X1 G5516 (
	 );
   AND3_X1 G5515 (
	 );
   NAND2_X1 G5514 (
	 );
   NAND2_X1 G5513 (
	 );
   NAND2_X1 G5512 (
	 );
   AOI22_X1 G5511 (
	 );
   AND3_X1 G5510 (
	 );
   NAND4_X1 G5509 (
	 );
   NAND4_X1 G5508 (
	 );
   NAND4_X1 G5507 (
	 );
   OAI21_X1 G5506 (
	 );
   INV_X1 G5505 (
	 );
   NAND2_X1 G5504 (
	 );
   CLKBUF_X1 G5503 (
	 );
   CLKBUF_X1 G5502 (
	 );
   NAND2_X1 G5501 (
	 );
   OAI21_X1 G5500 (
	 );
   NAND2_X1 G5499 (
	 );
   CLKBUF_X1 G5498 (
	 );
   OAI21_X1 G5497 (
	 );
   INV_X1 G5496 (
	 );
   CLKBUF_X1 G5495 (
	 );
   CLKBUF_X1 G5494 (
	 );
   CLKBUF_X1 G5493 (
	 );
   CLKBUF_X1 G5492 (
	 );
   CLKBUF_X1 G5491 (
	 );
   CLKBUF_X1 G5490 (
	 );
   CLKBUF_X1 G5489 (
	 );
   NAND4_X1 G5488 (
	 );
   NAND4_X1 G5487 (
	 );
   NAND4_X1 G5486 (
	 );
   NAND4_X1 G5485 (
	 );
   NOR2_X1 G5484 (
	 );
   AND2_X1 G5483 (
	 );
   NAND4_X1 G5482 (
	 );
   NAND4_X1 G5481 (
	 );
   NAND3_X1 G5480 (
	 );
   NAND3_X1 G5479 (
	 );
   NAND4_X1 G5478 (
	 );
   CLKBUF_X1 G5477 (
	 );
   CLKBUF_X1 G5476 (
	 );
   OAI21_X1 G5475 (
	 );
   INV_X1 G5474 (
	 );
   INV_X1 G5473 (
	 );
   NAND4_X1 G5472 (
	 );
   AOI22_X1 G5471 (
	 );
   NAND2_X1 G5470 (
	 );
   NAND2_X1 G5469 (
	 );
   NAND2_X1 G5468 (
	 );
   CLKBUF_X1 G5467 (
	 );
   OAI22_X1 G5466 (
	 );
   XNOR2_X1 G5465 (
	 );
   INV_X1 G5464 (
	 );
   CLKBUF_X1 G5463 (
	 );
   CLKBUF_X1 G5462 (
	 );
   CLKBUF_X1 G5461 (
	 );
   NOR3_X1 G5460 (
	 );
   AOI21_X1 G5459 (
	 );
   OAI21_X1 G5458 (
	 );
   NOR2_X1 G5457 (
	 );
   AND2_X1 G5456 (
	 );
   AOI21_X1 G5455 (
	 );
   INV_X1 G5454 (
	 );
   NOR2_X1 G5453 (
	 );
   CLKBUF_X1 G5452 (
	 );
   CLKBUF_X1 G5451 (
	 );
   CLKBUF_X1 G5450 (
	 );
   CLKBUF_X1 G5449 (
	 );
   AND2_X1 G5448 (
	 );
   OAI211_X1 G5447 (
	 );
   NOR2_X1 G5446 (
	 );
   NAND3_X1 G5445 (
	 );
   NAND4_X1 G5444 (
	 );
   OAI21_X1 G5443 (
	 );
   AOI21_X1 G5442 (
	 );
   OAI21_X1 G5441 (
	 );
   NOR2_X1 G5440 (
	 );
   AOI21_X1 G5439 (
	 );
   CLKBUF_X1 G5438 (
	 );
   CLKBUF_X1 G5437 (
	 );
   AOI221_X4 G5436 (
	 );
   NAND2_X1 G5435 (
	 );
   OAI21_X1 G5434 (
	 );
   NAND3_X1 G5433 (
	 );
   INV_X1 G5432 (
	 );
   NAND3_X1 G5431 (
	 );
   CLKBUF_X1 G5430 (
	 );
   MUX2_X1 G5429 (
	 );
   MUX2_X1 G5428 (
	 );
   CLKBUF_X1 G5427 (
	 );
   MUX2_X1 G5426 (
	 );
   OAI21_X1 G5425 (
	 );
   NAND2_X1 G5424 (
	 );
   MUX2_X1 G5423 (
	 );
   AND2_X1 G5422 (
	 );
   NOR2_X1 G5421 (
	 );
   CLKBUF_X1 G5420 (
	 );
   CLKBUF_X1 G5419 (
	 );
   OAI221_X1 G5418 (
	 );
   AOI22_X1 G5417 (
	 );
   CLKBUF_X1 G5416 (
	 );
   XNOR2_X1 G5415 (
	 );
   NAND2_X1 G5414 (
	 );
   CLKBUF_X1 G5413 (
	 );
   CLKBUF_X1 G5412 (
	 );
   NAND3_X1 G5411 (
	 );
   AOI22_X1 G5410 (
	 );
   AND3_X1 G5409 (
	 );
   NAND2_X1 G5408 (
	 );
   NAND2_X1 G5407 (
	 );
   NAND2_X1 G5406 (
	 );
   AND3_X1 G5405 (
	 );
   NAND4_X1 G5404 (
	 );
   NAND4_X1 G5403 (
	 );
   NAND4_X1 G5402 (
	 );
   NAND3_X1 G5401 (
	 );
   AOI22_X1 G5400 (
	 );
   AND3_X1 G5399 (
	 );
   NAND2_X1 G5398 (
	 );
   NAND2_X1 G5397 (
	 );
   NAND4_X1 G5396 (
	 );
   NAND3_X1 G5395 (
	 );
   NAND3_X1 G5394 (
	 );
   NAND3_X1 G5393 (
	 );
   NAND2_X1 G5392 (
	 );
   NAND2_X1 G5391 (
	 );
   AND3_X1 G5390 (
	 );
   NAND4_X1 G5389 (
	 );
   NAND4_X1 G5388 (
	 );
   NAND4_X1 G5387 (
	 );
   NOR4_X1 G5386 (
	 );
   CLKBUF_X1 G5385 (
	 );
   NOR2_X1 G5384 (
	 );
   XNOR2_X1 G5383 (
	 );
   NAND4_X1 G5382 (
	 );
   NAND3_X1 G5381 (
	 );
   NAND2_X1 G5380 (
	 );
   NAND2_X1 G5379 (
	 );
   OAI21_X1 G5378 (
	 );
   CLKBUF_X1 G5377 (
	 );
   CLKBUF_X1 G5376 (
	 );
   CLKBUF_X1 G5375 (
	 );
   MUX2_X1 G5374 (
	 );
   NOR3_X1 G5373 (
	 );
   INV_X1 G5372 (
	 );
   MUX2_X1 G5371 (
	 );
   CLKBUF_X1 G5370 (
	 );
   MUX2_X1 G5369 (
	 );
   CLKBUF_X1 G5368 (
	 );
   OAI21_X1 G5367 (
	 );
   INV_X1 G5366 (
	 );
   NAND2_X1 G5365 (
	 );
   CLKBUF_X1 G5364 (
	 );
   CLKBUF_X1 G5363 (
	 );
   CLKBUF_X1 G5362 (
	 );
   OAI21_X1 G5361 (
	 );
   INV_X1 G5360 (
	 );
   NAND2_X1 G5359 (
	 );
   OAI21_X1 G5358 (
	 );
   INV_X1 G5357 (
	 );
   NAND2_X1 G5356 (
	 );
   CLKBUF_X1 G5355 (
	 );
   CLKBUF_X1 G5354 (
	 );
   CLKBUF_X1 G5353 (
	 );
   NOR4_X1 G5352 (
	 );
   CLKBUF_X1 G5351 (
	 );
   CLKBUF_X1 G5350 (
	 );
   OAI21_X1 G5349 (
	 );
   INV_X1 G5348 (
	 );
   NAND2_X1 G5347 (
	 );
   NAND3_X1 G5346 (
	 );
   AOI22_X1 G5345 (
	 );
   AND3_X1 G5344 (
	 );
   NAND2_X1 G5343 (
	 );
   NAND2_X1 G5342 (
	 );
   NAND2_X1 G5341 (
	 );
   AND3_X1 G5340 (
	 );
   NAND4_X1 G5339 (
	 );
   NAND4_X1 G5338 (
	 );
   NAND4_X1 G5337 (
	 );
   CLKBUF_X1 G5336 (
	 );
   OAI21_X1 G5335 (
	 );
   NAND2_X1 G5334 (
	 );
   CLKBUF_X1 G5333 (
	 );
   AOI21_X1 G5332 (
	 );
   OAI21_X1 G5331 (
	 );
   NAND2_X1 G5330 (
	 );
   MUX2_X1 G5329 (
	 );
   NOR2_X1 G5328 (
	 );
   AOI21_X1 G5327 (
	 );
   NAND3_X1 G5326 (
	 );
   INV_X1 G5325 (
	 );
   AND2_X1 G5324 (
	 );
   OR4_X1 G5323 (
	 );
   NAND3_X1 G5322 (
	 );
   AOI22_X1 G5321 (
	 );
   AOI22_X1 G5320 (
	 );
   AOI22_X1 G5319 (
	 );
   NAND4_X1 G5318 (
	 );
   NAND2_X1 G5317 (
	 );
   AOI22_X1 G5316 (
	 );
   AOI22_X1 G5315 (
	 );
   AOI22_X1 G5314 (
	 );
   NAND4_X1 G5313 (
	 );
   AOI22_X1 G5312 (
	 );
   AOI22_X1 G5311 (
	 );
   AOI22_X1 G5310 (
	 );
   AOI22_X1 G5309 (
	 );
   NAND4_X1 G5308 (
	 );
   AOI22_X1 G5307 (
	 );
   AOI22_X1 G5306 (
	 );
   AOI22_X1 G5305 (
	 );
   AOI22_X1 G5304 (
	 );
   CLKBUF_X1 G5303 (
	 );
   CLKBUF_X1 G5302 (
	 );
   NAND2_X1 G5301 (
	 );
   AOI22_X1 G5300 (
	 );
   AOI22_X1 G5299 (
	 );
   CLKBUF_X1 G5298 (
	 );
   CLKBUF_X1 G5297 (
	 );
   CLKBUF_X1 G5296 (
	 );
   CLKBUF_X1 G5295 (
	 );
   MUX2_X1 G5294 (
	 );
   MUX2_X1 G5293 (
	 );
   CLKBUF_X1 G5292 (
	 );
   MUX2_X1 G5291 (
	 );
   OAI21_X1 G5290 (
	 );
   NAND2_X1 G5289 (
	 );
   OAI21_X1 G5288 (
	 );
   INV_X1 G5287 (
	 );
   NAND2_X1 G5286 (
	 );
   CLKBUF_X1 G5285 (
	 );
   NOR2_X1 G5284 (
	 );
   CLKBUF_X1 G5283 (
	 );
   CLKBUF_X1 G5282 (
	 );
   CLKBUF_X1 G5281 (
	 );
   CLKBUF_X1 G5280 (
	 );
   CLKBUF_X1 G5279 (
	 );
   OAI21_X1 G5278 (
	 );
   OAI21_X1 G5277 (
	 );
   NOR2_X1 G5276 (
	 );
   INV_X1 G5275 (
	 );
   NOR2_X1 G5274 (
	 );
   NAND2_X1 G5273 (
	 );
   AND2_X1 G5272 (
	 );
   CLKBUF_X1 G5271 (
	 );
   NAND4_X1 G5270 (
	 );
   NAND4_X1 G5269 (
	 );
   NAND4_X1 G5268 (
	 );
   NAND4_X1 G5267 (
	 );
   NOR2_X1 G5266 (
	 );
   NAND4_X1 G5265 (
	 );
   NAND4_X1 G5264 (
	 );
   NAND3_X1 G5263 (
	 );
   NAND3_X1 G5262 (
	 );
   NAND4_X1 G5261 (
	 );
   NAND2_X1 G5260 (
	 );
   NAND4_X1 G5259 (
	 );
   NAND4_X1 G5258 (
	 );
   AOI21_X1 G5257 (
	 );
   INV_X1 G5256 (
	 );
   CLKBUF_X1 G5255 (
	 );
   CLKBUF_X1 G5254 (
	 );
   CLKBUF_X1 G5253 (
	 );
   OAI21_X1 G5252 (
	 );
   INV_X1 G5251 (
	 );
   NAND2_X1 G5250 (
	 );
   OAI21_X1 G5249 (
	 );
   INV_X1 G5248 (
	 );
   NAND2_X1 G5247 (
	 );
   MUX2_X1 G5246 (
	 );
   CLKBUF_X1 G5245 (
	 );
   CLKBUF_X1 G5244 (
	 );
   CLKBUF_X1 G5243 (
	 );
   CLKBUF_X1 G5242 (
	 );
   CLKBUF_X1 G5241 (
	 );
   CLKBUF_X1 G5240 (
	 );
   CLKBUF_X1 G5239 (
	 );
   CLKBUF_X1 G5238 (
	 );
   CLKBUF_X1 G5237 (
	 );
   CLKBUF_X1 G5236 (
	 );
   CLKBUF_X1 G5235 (
	 );
   CLKBUF_X1 G5234 (
	 );
   CLKBUF_X1 G5233 (
	 );
   OAI21_X1 G5232 (
	 );
   NAND2_X1 G5231 (
	 );
   CLKBUF_X1 G5230 (
	 );
   CLKBUF_X1 G5229 (
	 );
   CLKBUF_X1 G5228 (
	 );
   AOI21_X1 G5227 (
	 );
   INV_X1 G5226 (
	 );
   NOR2_X1 G5225 (
	 );
   CLKBUF_X1 G5224 (
	 );
   NAND2_X1 G5223 (
	 );
   AOI22_X1 G5222 (
	 );
   AOI22_X1 G5221 (
	 );
   NOR2_X1 G5220 (
	 );
   AOI21_X1 G5219 (
	 );
   OAI21_X1 G5218 (
	 );
   NAND2_X1 G5217 (
	 );
   NOR2_X1 G5216 (
	 );
   AND2_X1 G5215 (
	 );
   CLKBUF_X1 G5214 (
	 );
   CLKBUF_X1 G5213 (
	 );
   CLKBUF_X1 G5212 (
	 );
   NAND3_X1 G5211 (
	 );
   AOI22_X1 G5210 (
	 );
   AND3_X1 G5209 (
	 );
   NAND2_X1 G5208 (
	 );
   NAND2_X1 G5207 (
	 );
   NAND2_X1 G5206 (
	 );
   AND3_X1 G5205 (
	 );
   NAND4_X1 G5204 (
	 );
   NAND4_X1 G5203 (
	 );
   NAND4_X1 G5202 (
	 );
   NAND2_X1 G5201 (
	 );
   NAND2_X1 G5200 (
	 );
   AOI22_X1 G5199 (
	 );
   NAND2_X1 G5198 (
	 );
   NAND3_X1 G5197 (
	 );
   OAI21_X1 G5196 (
	 );
   CLKBUF_X1 G5195 (
	 );
   OAI21_X1 G5194 (
	 );
   NAND2_X1 G5193 (
	 );
   OAI21_X1 G5192 (
	 );
   NOR2_X1 G5191 (
	 );
   CLKBUF_X1 G5190 (
	 );
   CLKBUF_X1 G5189 (
	 );
   CLKBUF_X1 G5188 (
	 );
   CLKBUF_X1 G5187 (
	 );
   CLKBUF_X1 G5186 (
	 );
   MUX2_X1 G5185 (
	 );
   NOR2_X1 G5184 (
	 );
   CLKBUF_X1 G5183 (
	 );
   NAND3_X1 G5182 (
	 );
   AOI22_X1 G5181 (
	 );
   AND3_X1 G5180 (
	 );
   NAND2_X1 G5179 (
	 );
   NAND2_X1 G5178 (
	 );
   NAND2_X1 G5177 (
	 );
   AND3_X1 G5176 (
	 );
   NAND4_X1 G5175 (
	 );
   NAND4_X1 G5174 (
	 );
   NAND4_X1 G5173 (
	 );
   NOR2_X1 G5172 (
	 );
   NOR2_X1 G5171 (
	 );
   NAND2_X1 G5170 (
	 );
   MUX2_X1 G5169 (
	 );
   AOI21_X1 G5168 (
	 );
   OAI21_X1 G5167 (
	 );
   CLKBUF_X1 G5166 (
	 );
   OAI221_X1 G5165 (
	 );
   AOI22_X1 G5164 (
	 );
   OAI21_X1 G5163 (
	 );
   INV_X1 G5162 (
	 );
   NAND2_X1 G5161 (
	 );
   CLKBUF_X1 G5160 (
	 );
   CLKBUF_X1 G5159 (
	 );
   AND2_X1 G5158 (
	 );
   CLKBUF_X1 G5157 (
	 );
   CLKBUF_X1 G5156 (
	 );
   CLKBUF_X1 G5155 (
	 );
   OAI21_X1 G5154 (
	 );
   INV_X1 G5153 (
	 );
   NAND2_X1 G5152 (
	 );
   OAI221_X1 G5151 (
	 );
   AOI22_X1 G5150 (
	 );
   CLKBUF_X1 G5149 (
	 );
   CLKBUF_X1 G5148 (
	 );
   CLKBUF_X1 G5147 (
	 );
   CLKBUF_X1 G5146 (
	 );
   MUX2_X1 G5145 (
	 );
   MUX2_X1 G5144 (
	 );
   CLKBUF_X1 G5143 (
	 );
   MUX2_X1 G5142 (
	 );
   CLKBUF_X1 G5141 (
	 );
   MUX2_X1 G5140 (
	 );
   MUX2_X1 G5139 (
	 );
   NAND2_X1 G5138 (
	 );
   AOI22_X1 G5137 (
	 );
   AOI22_X1 G5136 (
	 );
   CLKBUF_X1 G5135 (
	 );
   CLKBUF_X1 G5134 (
	 );
   CLKBUF_X1 G5133 (
	 );
   CLKBUF_X1 G5132 (
	 );
   MUX2_X1 G5131 (
	 );
   CLKBUF_X1 G5130 (
	 );
   CLKBUF_X1 G5129 (
	 );
   NOR2_X1 G5128 (
	 );
   CLKBUF_X1 G5127 (
	 );
   AOI21_X1 G5126 (
	 );
   INV_X1 G5125 (
	 );
   NOR2_X1 G5124 (
	 );
   CLKBUF_X1 G5123 (
	 );
   NAND2_X1 G5122 (
	 );
   AOI22_X1 G5121 (
	 );
   AOI22_X1 G5120 (
	 );
   CLKBUF_X1 G5119 (
	 );
   CLKBUF_X1 G5118 (
	 );
   OAI211_X1 G5117 (
	 );
   INV_X1 G5116 (
	 );
   NAND4_X1 G5115 (
	 );
   NOR3_X1 G5114 (
	 );
   AND3_X1 G5113 (
	 );
   NOR2_X1 G5112 (
	 );
   INV_X1 G5111 (
	 );
   OAI22_X1 G5110 (
	 );
   INV_X1 G5109 (
	 );
   INV_X1 G5108 (
	 );
   CLKBUF_X1 G5107 (
	 );
   CLKBUF_X1 G5106 (
	 );
   CLKBUF_X1 G5105 (
	 );
   CLKBUF_X1 G5104 (
	 );
   CLKBUF_X1 G5103 (
	 );
   OAI21_X1 G5102 (
	 );
   OR2_X1 G5101 (
	 );
   OAI211_X1 G5100 (
	 );
   OAI21_X1 G5099 (
	 );
   NAND2_X1 G5098 (
	 );
   MUX2_X1 G5097 (
	 );
   CLKBUF_X1 G5096 (
	 );
   MUX2_X1 G5095 (
	 );
   CLKBUF_X1 G5094 (
	 );
   OAI21_X1 G5093 (
	 );
   NAND2_X1 G5092 (
	 );
   CLKBUF_X1 G5091 (
	 );
   OAI221_X1 G5090 (
	 );
   AOI22_X1 G5089 (
	 );
   CLKBUF_X1 G5088 (
	 );
   CLKBUF_X1 G5087 (
	 );
   OAI21_X1 G5086 (
	 );
   INV_X1 G5085 (
	 );
   NAND2_X1 G5084 (
	 );
   OAI21_X1 G5083 (
	 );
   INV_X1 G5082 (
	 );
   NAND2_X1 G5081 (
	 );
   CLKBUF_X1 G5080 (
	 );
   CLKBUF_X1 G5079 (
	 );
   NOR2_X1 G5078 (
	 );
   CLKBUF_X1 G5077 (
	 );
   CLKBUF_X1 G5076 (
	 );
   NOR3_X1 G5075 (
	 );
   NOR2_X1 G5074 (
	 );
   NAND2_X1 G5073 (
	 );
   NAND2_X1 G5072 (
	 );
   AOI22_X1 G5071 (
	 );
   CLKBUF_X1 G5070 (
	 );
   CLKBUF_X1 G5069 (
	 );
   CLKBUF_X1 G5068 (
	 );
   NOR2_X1 G5067 (
	 );
   AND2_X1 G5066 (
	 );
   CLKBUF_X1 G5065 (
	 );
   CLKBUF_X1 G5064 (
	 );
   CLKBUF_X1 G5063 (
	 );
   CLKBUF_X1 G5062 (
	 );
   CLKBUF_X1 G5061 (
	 );
   AND2_X1 G5060 (
	 );
   CLKBUF_X1 G5059 (
	 );
   MUX2_X1 G5058 (
	 );
   OAI21_X1 G5057 (
	 );
   NAND2_X1 G5056 (
	 );
   OAI21_X1 G5055 (
	 );
   INV_X1 G5054 (
	 );
   INV_X1 G5053 (
	 );
   MUX2_X1 G5052 (
	 );
   CLKBUF_X1 G5051 (
	 );
   OAI221_X1 G5050 (
	 );
   AOI22_X1 G5049 (
	 );
   CLKBUF_X1 G5048 (
	 );
   CLKBUF_X1 G5047 (
	 );
   OAI21_X1 G5046 (
	 );
   INV_X1 G5045 (
	 );
   NAND2_X1 G5044 (
	 );
   CLKBUF_X1 G5043 (
	 );
   NAND4_X1 G5042 (
	 );
   INV_X1 G5041 (
	 );
   CLKBUF_X1 G5040 (
	 );
   CLKBUF_X1 G5039 (
	 );
   CLKBUF_X1 G5038 (
	 );
   CLKBUF_X1 G5037 (
	 );
   CLKBUF_X1 G5036 (
	 );
   CLKBUF_X1 G5035 (
	 );
   OAI21_X1 G5034 (
	 );
   INV_X1 G5033 (
	 );
   NAND2_X1 G5032 (
	 );
   OAI22_X1 G5031 (
	 );
   XNOR2_X1 G5030 (
	 );
   INV_X1 G5029 (
	 );
   NOR2_X1 G5028 (
	 );
   AOI21_X1 G5027 (
	 );
   NAND2_X1 G5026 (
	 );
   NAND2_X1 G5025 (
	 );
   OAI211_X1 G5024 (
	 );
   CLKBUF_X1 G5023 (
	 );
   AND2_X1 G5022 (
	 );
   CLKBUF_X1 G5021 (
	 );
   MUX2_X1 G5020 (
	 );
   OAI21_X1 G5019 (
	 );
   NAND2_X1 G5018 (
	 );
   MUX2_X1 G5017 (
	 );
   CLKBUF_X1 G5016 (
	 );
   AND2_X1 G5015 (
	 );
   NAND4_X1 G5014 (
	 );
   NAND2_X1 G5013 (
	 );
   AOI22_X1 G5012 (
	 );
   NAND2_X1 G5011 (
	 );
   NAND2_X1 G5010 (
	 );
   OAI211_X1 G5009 (
	 );
   NAND3_X1 G5008 (
	 );
   OAI21_X1 G5007 (
	 );
   OAI21_X1 G5006 (
	 );
   NAND2_X1 G5005 (
	 );
   CLKBUF_X1 G5004 (
	 );
   NOR2_X1 G5003 (
	 );
   NAND3_X1 G5002 (
	 );
   OR2_X1 G5001 (
	 );
   NOR3_X1 G5000 (
	 );
   NAND3_X1 G4999 (
	 );
   NAND4_X1 G4998 (
	 );
   NAND3_X1 G4997 (
	 );
   NAND3_X1 G4996 (
	 );
   OAI22_X1 G4995 (
	 );
   INV_X1 G4994 (
	 );
   AND4_X1 G4993 (
	 );
   NOR2_X1 G4992 (
	 );
   NOR2_X1 G4991 (
	 );
   NOR2_X1 G4990 (
	 );
   INV_X1 G4989 (
	 );
   MUX2_X1 G4988 (
	 );
   CLKBUF_X1 G4987 (
	 );
   OAI21_X1 G4986 (
	 );
   INV_X1 G4985 (
	 );
   NAND2_X1 G4984 (
	 );
   MUX2_X1 G4983 (
	 );
   CLKBUF_X1 G4982 (
	 );
   CLKBUF_X1 G4981 (
	 );
   NOR2_X1 G4980 (
	 );
   OAI21_X1 G4979 (
	 );
   INV_X1 G4978 (
	 );
   NAND2_X1 G4977 (
	 );
   NOR2_X1 G4976 (
	 );
   OAI221_X1 G4975 (
	 );
   AOI22_X1 G4974 (
	 );
   CLKBUF_X1 G4973 (
	 );
   CLKBUF_X1 G4972 (
	 );
   CLKBUF_X1 G4971 (
	 );
   NAND3_X1 G4970 (
	 );
   AOI22_X1 G4969 (
	 );
   AND3_X1 G4968 (
	 );
   NAND2_X1 G4967 (
	 );
   NAND2_X1 G4966 (
	 );
   NAND2_X1 G4965 (
	 );
   AND3_X1 G4964 (
	 );
   NAND4_X1 G4963 (
	 );
   NAND4_X1 G4962 (
	 );
   NAND4_X1 G4961 (
	 );
   CLKBUF_X1 G4960 (
	 );
   CLKBUF_X1 G4959 (
	 );
   CLKBUF_X1 G4958 (
	 );
   CLKBUF_X1 G4957 (
	 );
   AOI21_X1 G4956 (
	 );
   NOR2_X1 G4955 (
	 );
   CLKBUF_X1 G4954 (
	 );
   NOR2_X1 G4953 (
	 );
   INV_X1 G4952 (
	 );
   CLKBUF_X1 G4951 (
	 );
   OAI221_X1 G4950 (
	 );
   INV_X1 G4949 (
	 );
   INV_X1 G4948 (
	 );
   AOI22_X1 G4947 (
	 );
   OAI21_X1 G4946 (
	 );
   INV_X1 G4945 (
	 );
   NAND2_X1 G4944 (
	 );
   CLKBUF_X1 G4943 (
	 );
   MUX2_X1 G4942 (
	 );
   NOR2_X1 G4941 (
	 );
   NAND2_X1 G4940 (
	 );
   AND2_X1 G4939 (
	 );
   CLKBUF_X1 G4938 (
	 );
   CLKBUF_X1 G4937 (
	 );
   MUX2_X1 G4936 (
	 );
   CLKBUF_X1 G4935 (
	 );
   CLKBUF_X1 G4934 (
	 );
   OAI221_X1 G4933 (
	 );
   INV_X1 G4932 (
	 );
   AOI22_X1 G4931 (
	 );
   CLKBUF_X1 G4930 (
	 );
   CLKBUF_X1 G4929 (
	 );
   CLKBUF_X1 G4928 (
	 );
   NAND2_X1 G4927 (
	 );
   AOI22_X1 G4926 (
	 );
   AOI22_X1 G4925 (
	 );
   CLKBUF_X1 G4924 (
	 );
   OAI21_X1 G4923 (
	 );
   NAND2_X1 G4922 (
	 );
   OAI21_X1 G4921 (
	 );
   NAND2_X1 G4920 (
	 );
   CLKBUF_X1 G4919 (
	 );
   MUX2_X1 G4918 (
	 );
   CLKBUF_X1 G4917 (
	 );
   NOR3_X1 G4916 (
	 );
   AOI21_X1 G4915 (
	 );
   CLKBUF_X1 G4914 (
	 );
   MUX2_X1 G4913 (
	 );
   CLKBUF_X1 G4912 (
	 );
   CLKBUF_X1 G4911 (
	 );
   NAND3_X1 G4910 (
	 );
   AOI22_X1 G4909 (
	 );
   NAND4_X1 G4908 (
	 );
   NAND3_X1 G4907 (
	 );
   NAND3_X1 G4906 (
	 );
   NAND3_X1 G4905 (
	 );
   NAND2_X1 G4904 (
	 );
   AND3_X1 G4903 (
	 );
   NAND2_X1 G4902 (
	 );
   NAND2_X1 G4901 (
	 );
   NAND2_X1 G4900 (
	 );
   AND3_X1 G4899 (
	 );
   NAND4_X1 G4898 (
	 );
   NAND4_X1 G4897 (
	 );
   NAND4_X1 G4896 (
	 );
   OAI21_X1 G4895 (
	 );
   INV_X1 G4894 (
	 );
   NAND2_X1 G4893 (
	 );
   CLKBUF_X1 G4892 (
	 );
   CLKBUF_X1 G4891 (
	 );
   CLKBUF_X1 G4890 (
	 );
   CLKBUF_X1 G4889 (
	 );
   CLKBUF_X1 G4888 (
	 );
   NOR2_X1 G4887 (
	 );
   AND2_X1 G4886 (
	 );
   NOR3_X1 G4885 (
	 );
   CLKBUF_X1 G4884 (
	 );
   NAND4_X1 G4883 (
	 );
   NAND4_X1 G4882 (
	 );
   OR2_X1 G4881 (
	 );
   OR2_X1 G4880 (
	 );
   NOR2_X1 G4879 (
	 );
   AND2_X1 G4878 (
	 );
   NAND4_X1 G4877 (
	 );
   NAND4_X1 G4876 (
	 );
   NAND3_X1 G4875 (
	 );
   NAND3_X1 G4874 (
	 );
   NAND4_X1 G4873 (
	 );
   CLKBUF_X1 G4872 (
	 );
   NAND4_X1 G4871 (
	 );
   NAND2_X1 G4870 (
	 );
   NAND2_X1 G4869 (
	 );
   NAND2_X1 G4868 (
	 );
   AOI22_X1 G4867 (
	 );
   CLKBUF_X1 G4866 (
	 );
   CLKBUF_X1 G4865 (
	 );
   CLKBUF_X1 G4864 (
	 );
   OAI21_X1 G4863 (
	 );
   INV_X1 G4862 (
	 );
   NAND2_X1 G4861 (
	 );
   NOR2_X1 G4860 (
	 );
   NOR3_X1 G4859 (
	 );
   NOR3_X1 G4858 (
	 );
   CLKBUF_X1 G4857 (
	 );
   MUX2_X1 G4856 (
	 );
   CLKBUF_X1 G4855 (
	 );
   OAI21_X1 G4854 (
	 );
   NAND2_X1 G4853 (
	 );
   OAI21_X1 G4852 (
	 );
   NOR2_X1 G4851 (
	 );
   NOR2_X1 G4850 (
	 );
   MUX2_X1 G4849 (
	 );
   AOI21_X1 G4848 (
	 );
   INV_X1 G4847 (
	 );
   OAI221_X1 G4846 (
	 );
   NAND2_X1 G4845 (
	 );
   OAI21_X1 G4844 (
	 );
   NAND3_X1 G4843 (
	 );
   XOR2_X1 G4842 (
	 );
   NOR2_X1 G4841 (
	 );
   AND2_X1 G4840 (
	 );
   CLKBUF_X1 G4839 (
	 );
   NOR2_X1 G4838 (
	 );
   NOR3_X1 G4837 (
	 );
   NOR3_X1 G4836 (
	 );
   CLKBUF_X1 G4835 (
	 );
   NAND2_X1 G4834 (
	 );
   AND4_X1 G4833 (
	 );
   NAND2_X1 G4832 (
	 );
   NAND2_X1 G4831 (
	 );
   NAND4_X1 G4830 (
	 );
   NAND3_X1 G4829 (
	 );
   NAND3_X1 G4828 (
	 );
   NAND3_X1 G4827 (
	 );
   NAND2_X1 G4826 (
	 );
   NAND2_X1 G4825 (
	 );
   NAND2_X1 G4824 (
	 );
   AND4_X1 G4823 (
	 );
   NAND4_X1 G4822 (
	 );
   NAND4_X1 G4821 (
	 );
   NAND3_X1 G4820 (
	 );
   NAND3_X1 G4819 (
	 );
   CLKBUF_X1 G4818 (
	 );
   CLKBUF_X1 G4817 (
	 );
   CLKBUF_X1 G4816 (
	 );
   CLKBUF_X1 G4815 (
	 );
   AND2_X1 G4814 (
	 );
   CLKBUF_X1 G4813 (
	 );
   CLKBUF_X1 G4812 (
	 );
   CLKBUF_X1 G4811 (
	 );
   CLKBUF_X1 G4810 (
	 );
   CLKBUF_X1 G4809 (
	 );
   MUX2_X1 G4808 (
	 );
   MUX2_X1 G4807 (
	 );
   CLKBUF_X1 G4806 (
	 );
   OAI22_X1 G4805 (
	 );
   INV_X1 G4804 (
	 );
   XNOR2_X1 G4803 (
	 );
   CLKBUF_X1 G4802 (
	 );
   CLKBUF_X1 G4801 (
	 );
   CLKBUF_X1 G4800 (
	 );
   CLKBUF_X1 G4799 (
	 );
   NOR2_X1 G4798 (
	 );
   OAI221_X1 G4797 (
	 );
   AOI22_X1 G4796 (
	 );
   AOI21_X1 G4795 (
	 );
   INV_X1 G4794 (
	 );
   NOR2_X1 G4793 (
	 );
   CLKBUF_X1 G4792 (
	 );
   CLKBUF_X1 G4791 (
	 );
   CLKBUF_X1 G4790 (
	 );
   MUX2_X1 G4789 (
	 );
   CLKBUF_X1 G4788 (
	 );
   CLKBUF_X1 G4787 (
	 );
   INV_X1 G4786 (
	 );
   CLKBUF_X1 G4785 (
	 );
   MUX2_X1 G4784 (
	 );
   AND2_X1 G4783 (
	 );
   INV_X1 G4782 (
	 );
   AOI211_X1 G4781 (
	 );
   CLKBUF_X1 G4780 (
	 );
   NAND3_X1 G4779 (
	 );
   AOI22_X1 G4778 (
	 );
   AND3_X1 G4777 (
	 );
   NAND2_X1 G4776 (
	 );
   NAND2_X1 G4775 (
	 );
   NAND2_X1 G4774 (
	 );
   AND3_X1 G4773 (
	 );
   NAND4_X1 G4772 (
	 );
   NAND4_X1 G4771 (
	 );
   NAND4_X1 G4770 (
	 );
   AOI21_X1 G4769 (
	 );
   INV_X1 G4768 (
	 );
   NOR2_X1 G4767 (
	 );
   CLKBUF_X1 G4766 (
	 );
   CLKBUF_X1 G4765 (
	 );
   OAI221_X1 G4764 (
	 );
   INV_X1 G4763 (
	 );
   INV_X1 G4762 (
	 );
   AOI22_X1 G4761 (
	 );
   CLKBUF_X1 G4760 (
	 );
   NAND2_X1 G4759 (
	 );
   AOI22_X1 G4758 (
	 );
   AOI22_X1 G4757 (
	 );
   CLKBUF_X1 G4756 (
	 );
   NAND2_X1 G4755 (
	 );
   AOI22_X1 G4754 (
	 );
   AOI22_X1 G4753 (
	 );
   NOR2_X1 G4752 (
	 );
   NOR2_X1 G4751 (
	 );
   NAND3_X1 G4750 (
	 );
   CLKBUF_X1 G4749 (
	 );
   CLKBUF_X1 G4748 (
	 );
   CLKBUF_X1 G4747 (
	 );
   MUX2_X1 G4746 (
	 );
   OAI21_X1 G4745 (
	 );
   NAND2_X1 G4744 (
	 );
   CLKBUF_X1 G4743 (
	 );
   MUX2_X1 G4742 (
	 );
   CLKBUF_X1 G4741 (
	 );
   NAND2_X1 G4740 (
	 );
   AND4_X1 G4739 (
	 );
   NAND2_X1 G4738 (
	 );
   NAND2_X1 G4737 (
	 );
   NAND2_X1 G4736 (
	 );
   NAND2_X1 G4735 (
	 );
   AND4_X1 G4734 (
	 );
   NAND4_X1 G4733 (
	 );
   NAND4_X1 G4732 (
	 );
   NAND3_X1 G4731 (
	 );
   NAND3_X1 G4730 (
	 );
   OAI21_X1 G4729 (
	 );
   INV_X1 G4728 (
	 );
   NAND2_X1 G4727 (
	 );
   OAI21_X1 G4726 (
	 );
   INV_X1 G4725 (
	 );
   NAND2_X1 G4724 (
	 );
   MUX2_X1 G4723 (
	 );
   CLKBUF_X1 G4722 (
	 );
   CLKBUF_X1 G4721 (
	 );
   CLKBUF_X1 G4720 (
	 );
   OAI21_X1 G4719 (
	 );
   INV_X1 G4718 (
	 );
   NAND2_X1 G4717 (
	 );
   CLKBUF_X1 G4716 (
	 );
   CLKBUF_X1 G4715 (
	 );
   CLKBUF_X1 G4714 (
	 );
   CLKBUF_X1 G4713 (
	 );
   CLKBUF_X1 G4712 (
	 );
   CLKBUF_X1 G4711 (
	 );
   CLKBUF_X1 G4710 (
	 );
   CLKBUF_X1 G4709 (
	 );
   NAND2_X1 G4708 (
	 );
   NOR2_X1 G4707 (
	 );
   NAND3_X1 G4706 (
	 );
   AND3_X1 G4705 (
	 );
   NAND2_X1 G4704 (
	 );
   NAND2_X1 G4703 (
	 );
   NAND2_X1 G4702 (
	 );
   AOI22_X1 G4701 (
	 );
   AND3_X1 G4700 (
	 );
   NAND4_X1 G4699 (
	 );
   NAND4_X1 G4698 (
	 );
   NAND4_X1 G4697 (
	 );
   CLKBUF_X1 G4696 (
	 );
   AND2_X1 G4695 (
	 );
   MUX2_X1 G4694 (
	 );
   CLKBUF_X1 G4693 (
	 );
   AOI21_X1 G4692 (
	 );
   INV_X1 G4691 (
	 );
   NAND3_X1 G4690 (
	 );
   AOI21_X1 G4689 (
	 );
   AOI21_X1 G4688 (
	 );
   OAI21_X1 G4687 (
	 );
   INV_X1 G4686 (
	 );
   NOR2_X1 G4685 (
	 );
   CLKBUF_X1 G4684 (
	 );
   CLKBUF_X1 G4683 (
	 );
   CLKBUF_X1 G4682 (
	 );
   CLKBUF_X1 G4681 (
	 );
   CLKBUF_X1 G4680 (
	 );
   AOI21_X1 G4679 (
	 );
   INV_X1 G4678 (
	 );
   NOR2_X1 G4677 (
	 );
   OAI221_X1 G4676 (
	 );
   INV_X1 G4675 (
	 );
   INV_X1 G4674 (
	 );
   AOI22_X1 G4673 (
	 );
   NOR2_X1 G4672 (
	 );
   AOI21_X1 G4671 (
	 );
   NOR2_X1 G4670 (
	 );
   CLKBUF_X1 G4669 (
	 );
   CLKBUF_X1 G4668 (
	 );
   CLKBUF_X1 G4667 (
	 );
   CLKBUF_X1 G4666 (
	 );
   AOI21_X1 G4665 (
	 );
   NAND3_X1 G4664 (
	 );
   INV_X1 G4663 (
	 );
   CLKBUF_X1 G4662 (
	 );
   CLKBUF_X1 G4661 (
	 );
   CLKBUF_X1 G4660 (
	 );
   NAND2_X1 G4659 (
	 );
   AOI22_X1 G4658 (
	 );
   AOI22_X1 G4657 (
	 );
   CLKBUF_X1 G4656 (
	 );
   NOR2_X1 G4655 (
	 );
   CLKBUF_X1 G4654 (
	 );
   CLKBUF_X1 G4653 (
	 );
   AOI21_X1 G4652 (
	 );
   OAI21_X1 G4651 (
	 );
   NAND2_X1 G4650 (
	 );
   CLKBUF_X1 G4649 (
	 );
   MUX2_X1 G4648 (
	 );
   NOR2_X1 G4647 (
	 );
   AOI21_X1 G4646 (
	 );
   CLKBUF_X1 G4645 (
	 );
   OAI21_X1 G4644 (
	 );
   NAND2_X1 G4643 (
	 );
   CLKBUF_X1 G4642 (
	 );
   AND2_X1 G4641 (
	 );
   CLKBUF_X1 G4640 (
	 );
   CLKBUF_X1 G4639 (
	 );
   CLKBUF_X1 G4638 (
	 );
   OAI21_X1 G4637 (
	 );
   NOR2_X1 G4636 (
	 );
   NOR2_X1 G4635 (
	 );
   OAI221_X1 G4634 (
	 );
   INV_X1 G4633 (
	 );
   AOI22_X1 G4632 (
	 );
   CLKBUF_X1 G4631 (
	 );
   OAI211_X1 G4630 (
	 );
   NAND4_X1 G4629 (
	 );
   NOR3_X1 G4628 (
	 );
   AND3_X1 G4627 (
	 );
   NOR2_X1 G4626 (
	 );
   INV_X1 G4625 (
	 );
   OAI22_X1 G4624 (
	 );
   INV_X1 G4623 (
	 );
   INV_X1 G4622 (
	 );
   CLKBUF_X1 G4621 (
	 );
   AOI21_X1 G4620 (
	 );
   INV_X1 G4619 (
	 );
   NOR2_X1 G4618 (
	 );
   CLKBUF_X1 G4617 (
	 );
   CLKBUF_X1 G4616 (
	 );
   XNOR2_X1 G4615 (
	 );
   NAND2_X1 G4614 (
	 );
   XNOR2_X1 G4613 (
	 );
   CLKBUF_X1 G4612 (
	 );
   CLKBUF_X1 G4611 (
	 );
   CLKBUF_X1 G4610 (
	 );
   CLKBUF_X1 G4609 (
	 );
   CLKBUF_X1 G4608 (
	 );
   OAI21_X1 G4607 (
	 );
   INV_X1 G4606 (
	 );
   NAND2_X1 G4605 (
	 );
   OAI21_X1 G4604 (
	 );
   NAND2_X1 G4603 (
	 );
   NAND2_X1 G4602 (
	 );
   INV_X1 G4601 (
	 );
   NAND3_X1 G4600 (
	 );
   AOI22_X1 G4599 (
	 );
   AND3_X1 G4598 (
	 );
   NAND2_X1 G4597 (
	 );
   NAND2_X1 G4596 (
	 );
   NAND2_X1 G4595 (
	 );
   AND3_X1 G4594 (
	 );
   NAND4_X1 G4593 (
	 );
   NAND4_X1 G4592 (
	 );
   NAND4_X1 G4591 (
	 );
   CLKBUF_X1 G4590 (
	 );
   CLKBUF_X1 G4589 (
	 );
   CLKBUF_X1 G4588 (
	 );
   NAND4_X1 G4587 (
	 );
   NAND4_X1 G4586 (
	 );
   OR2_X1 G4585 (
	 );
   OR2_X1 G4584 (
	 );
   NOR2_X1 G4583 (
	 );
   NOR2_X1 G4582 (
	 );
   NAND4_X1 G4581 (
	 );
   NAND4_X1 G4580 (
	 );
   NAND3_X1 G4579 (
	 );
   NAND3_X1 G4578 (
	 );
   NAND4_X1 G4577 (
	 );
   MUX2_X1 G4576 (
	 );
   CLKBUF_X1 G4575 (
	 );
   CLKBUF_X1 G4574 (
	 );
   CLKBUF_X1 G4573 (
	 );
   MUX2_X1 G4572 (
	 );
   AOI21_X1 G4571 (
	 );
   OAI21_X1 G4570 (
	 );
   NOR4_X1 G4569 (
	 );
   NAND3_X1 G4568 (
	 );
   NAND4_X1 G4567 (
	 );
   NOR3_X1 G4566 (
	 );
   NAND3_X1 G4565 (
	 );
   NAND4_X1 G4564 (
	 );
   NAND3_X1 G4563 (
	 );
   NAND3_X1 G4562 (
	 );
   OAI22_X1 G4561 (
	 );
   INV_X1 G4560 (
	 );
   AND4_X1 G4559 (
	 );
   NOR2_X1 G4558 (
	 );
   NOR2_X1 G4557 (
	 );
   INV_X1 G4556 (
	 );
   NOR2_X1 G4555 (
	 );
   INV_X1 G4554 (
	 );
   AND2_X1 G4553 (
	 );
   OAI21_X1 G4552 (
	 );
   NAND2_X1 G4551 (
	 );
   AOI21_X1 G4550 (
	 );
   INV_X1 G4549 (
	 );
   NOR2_X1 G4548 (
	 );
   CLKBUF_X1 G4547 (
	 );
   CLKBUF_X1 G4546 (
	 );
   AOI21_X1 G4545 (
	 );
   CLKBUF_X1 G4544 (
	 );
   CLKBUF_X1 G4543 (
	 );
   MUX2_X1 G4542 (
	 );
   NAND2_X1 G4541 (
	 );
   AOI22_X1 G4540 (
	 );
   AOI22_X1 G4539 (
	 );
   MUX2_X1 G4538 (
	 );
   NAND3_X1 G4537 (
	 );
   AOI22_X1 G4536 (
	 );
   AND3_X1 G4535 (
	 );
   NAND2_X1 G4534 (
	 );
   NAND2_X1 G4533 (
	 );
   NAND2_X1 G4532 (
	 );
   AND3_X1 G4531 (
	 );
   NAND4_X1 G4530 (
	 );
   NAND4_X1 G4529 (
	 );
   NAND4_X1 G4528 (
	 );
   NAND4_X1 G4527 (
	 );
   AOI22_X1 G4526 (
	 );
   NAND2_X1 G4525 (
	 );
   NAND4_X1 G4524 (
	 );
   NAND3_X1 G4523 (
	 );
   NAND3_X1 G4522 (
	 );
   NAND3_X1 G4521 (
	 );
   NAND2_X1 G4520 (
	 );
   NAND2_X1 G4519 (
	 );
   NAND2_X1 G4518 (
	 );
   AOI22_X1 G4517 (
	 );
   AOI22_X1 G4516 (
	 );
   NAND2_X1 G4515 (
	 );
   AOI21_X1 G4514 (
	 );
   NOR2_X1 G4513 (
	 );
   INV_X1 G4512 (
	 );
   NOR3_X1 G4511 (
	 );
   NOR2_X1 G4510 (
	 );
   CLKBUF_X1 G4509 (
	 );
   CLKBUF_X1 G4508 (
	 );
   AND2_X1 G4507 (
	 );
   CLKBUF_X1 G4506 (
	 );
   MUX2_X1 G4505 (
	 );
   AND2_X1 G4504 (
	 );
   OAI21_X1 G4503 (
	 );
   INV_X1 G4502 (
	 );
   NAND2_X1 G4501 (
	 );
   NOR2_X1 G4500 (
	 );
   AND2_X1 G4499 (
	 );
   CLKBUF_X1 G4498 (
	 );
   OAI221_X1 G4497 (
	 );
   AOI22_X1 G4496 (
	 );
   OAI221_X1 G4495 (
	 );
   OAI21_X1 G4494 (
	 );
   CLKBUF_X1 G4493 (
	 );
   AND2_X1 G4492 (
	 );
   OAI221_X1 G4491 (
	 );
   INV_X1 G4490 (
	 );
   AOI22_X1 G4489 (
	 );
   MUX2_X1 G4488 (
	 );
   MUX2_X1 G4487 (
	 );
   CLKBUF_X1 G4486 (
	 );
   CLKBUF_X1 G4485 (
	 );
   NAND2_X1 G4484 (
	 );
   NAND2_X1 G4483 (
	 );
   AOI22_X1 G4482 (
	 );
   CLKBUF_X1 G4481 (
	 );
   OAI21_X1 G4480 (
	 );
   NAND2_X1 G4479 (
	 );
   AOI21_X1 G4478 (
	 );
   AOI21_X1 G4477 (
	 );
   NAND2_X1 G4476 (
	 );
   AOI21_X1 G4475 (
	 );
   NOR2_X1 G4474 (
	 );
   CLKBUF_X1 G4473 (
	 );
   NAND2_X1 G4472 (
	 );
   AOI22_X1 G4471 (
	 );
   AOI22_X1 G4470 (
	 );
   OAI221_X1 G4469 (
	 );
   INV_X1 G4468 (
	 );
   INV_X1 G4467 (
	 );
   AOI22_X1 G4466 (
	 );
   NAND3_X1 G4465 (
	 );
   NAND4_X1 G4464 (
	 );
   NOR3_X1 G4463 (
	 );
   NAND3_X1 G4462 (
	 );
   NAND4_X1 G4461 (
	 );
   NAND3_X1 G4460 (
	 );
   NAND3_X1 G4459 (
	 );
   OAI22_X1 G4458 (
	 );
   INV_X1 G4457 (
	 );
   AND4_X1 G4456 (
	 );
   NOR2_X1 G4455 (
	 );
   NOR2_X1 G4454 (
	 );
   INV_X1 G4453 (
	 );
   NOR2_X1 G4452 (
	 );
   INV_X1 G4451 (
	 );
   CLKBUF_X1 G4450 (
	 );
   CLKBUF_X1 G4449 (
	 );
   CLKBUF_X1 G4448 (
	 );
   CLKBUF_X1 G4447 (
	 );
   OAI21_X1 G4446 (
	 );
   INV_X1 G4445 (
	 );
   NAND2_X1 G4444 (
	 );
   CLKBUF_X1 G4443 (
	 );
   CLKBUF_X1 G4442 (
	 );
   CLKBUF_X1 G4441 (
	 );
   NOR2_X1 G4440 (
	 );
   NAND4_X1 G4439 (
	 );
   NAND2_X1 G4438 (
	 );
   NAND2_X1 G4437 (
	 );
   NAND2_X1 G4436 (
	 );
   AOI22_X1 G4435 (
	 );
   CLKBUF_X1 G4434 (
	 );
   NOR3_X1 G4433 (
	 );
   AOI21_X1 G4432 (
	 );
   CLKBUF_X1 G4431 (
	 );
   OAI21_X1 G4430 (
	 );
   NAND2_X1 G4429 (
	 );
   AND2_X1 G4428 (
	 );
   CLKBUF_X1 G4427 (
	 );
   CLKBUF_X1 G4426 (
	 );
   OAI21_X1 G4425 (
	 );
   INV_X1 G4424 (
	 );
   NAND2_X1 G4423 (
	 );
   MUX2_X1 G4422 (
	 );
   CLKBUF_X1 G4421 (
	 );
   CLKBUF_X1 G4420 (
	 );
   CLKBUF_X1 G4419 (
	 );
   NAND4_X1 G4418 (
	 );
   NAND2_X1 G4417 (
	 );
   NAND2_X1 G4416 (
	 );
   NAND2_X1 G4415 (
	 );
   AOI22_X1 G4414 (
	 );
   INV_X1 G4413 (
	 );
   CLKBUF_X1 G4412 (
	 );
   AOI21_X1 G4411 (
	 );
   OAI21_X1 G4410 (
	 );
   NAND2_X1 G4409 (
	 );
   CLKBUF_X1 G4408 (
	 );
   CLKBUF_X1 G4407 (
	 );
   CLKBUF_X1 G4406 (
	 );
   CLKBUF_X1 G4405 (
	 );
   OAI21_X1 G4404 (
	 );
   NAND2_X1 G4403 (
	 );
   MUX2_X1 G4402 (
	 );
   CLKBUF_X1 G4401 (
	 );
   OAI21_X1 G4400 (
	 );
   INV_X1 G4399 (
	 );
   NAND2_X1 G4398 (
	 );
   MUX2_X1 G4397 (
	 );
   CLKBUF_X1 G4396 (
	 );
   CLKBUF_X1 G4395 (
	 );
   CLKBUF_X1 G4394 (
	 );
   OAI221_X1 G4393 (
	 );
   INV_X1 G4392 (
	 );
   INV_X1 G4391 (
	 );
   AOI22_X1 G4390 (
	 );
   CLKBUF_X1 G4389 (
	 );
   NAND2_X1 G4388 (
	 );
   AOI22_X1 G4387 (
	 );
   AOI22_X1 G4386 (
	 );
   CLKBUF_X1 G4385 (
	 );
   CLKBUF_X1 G4384 (
	 );
   NAND3_X1 G4383 (
	 );
   AOI22_X1 G4382 (
	 );
   AND3_X1 G4381 (
	 );
   NAND2_X1 G4380 (
	 );
   NAND2_X1 G4379 (
	 );
   NAND2_X1 G4378 (
	 );
   AND3_X1 G4377 (
	 );
   NAND4_X1 G4376 (
	 );
   NAND4_X1 G4375 (
	 );
   NAND4_X1 G4374 (
	 );
   CLKBUF_X1 G4373 (
	 );
   CLKBUF_X1 G4372 (
	 );
   CLKBUF_X1 G4371 (
	 );
   OAI21_X1 G4370 (
	 );
   NAND2_X1 G4369 (
	 );
   CLKBUF_X1 G4368 (
	 );
   CLKBUF_X1 G4367 (
	 );
   MUX2_X1 G4366 (
	 );
   AND2_X1 G4365 (
	 );
   MUX2_X1 G4364 (
	 );
   CLKBUF_X1 G4363 (
	 );
   CLKBUF_X1 G4362 (
	 );
   CLKBUF_X1 G4361 (
	 );
   NAND2_X1 G4360 (
	 );
   NAND2_X1 G4359 (
	 );
   AND2_X1 G4358 (
	 );
   NAND4_X1 G4357 (
	 );
   AOI22_X1 G4356 (
	 );
   NAND2_X1 G4355 (
	 );
   NAND2_X1 G4354 (
	 );
   NAND2_X1 G4353 (
	 );
   CLKBUF_X1 G4352 (
	 );
   CLKBUF_X1 G4351 (
	 );
   CLKBUF_X1 G4350 (
	 );
   CLKBUF_X1 G4349 (
	 );
   OAI22_X1 G4348 (
	 );
   NAND2_X1 G4347 (
	 );
   INV_X1 G4346 (
	 );
   OAI21_X1 G4345 (
	 );
   INV_X1 G4344 (
	 );
   NAND2_X1 G4343 (
	 );
   AND2_X1 G4342 (
	 );
   CLKBUF_X1 G4341 (
	 );
   AND2_X1 G4340 (
	 );
   AND2_X1 G4339 (
	 );
   OAI21_X1 G4338 (
	 );
   NAND2_X1 G4337 (
	 );
   CLKBUF_X1 G4336 (
	 );
   NAND3_X1 G4335 (
	 );
   AND3_X1 G4334 (
	 );
   NAND2_X1 G4333 (
	 );
   NAND2_X1 G4332 (
	 );
   NAND2_X1 G4331 (
	 );
   AOI22_X1 G4330 (
	 );
   AND3_X1 G4329 (
	 );
   NAND4_X1 G4328 (
	 );
   NAND4_X1 G4327 (
	 );
   NAND4_X1 G4326 (
	 );
   CLKBUF_X1 G4325 (
	 );
   CLKBUF_X1 G4324 (
	 );
   OAI221_X1 G4323 (
	 );
   OAI21_X1 G4322 (
	 );
   CLKBUF_X1 G4321 (
	 );
   NOR2_X1 G4320 (
	 );
   CLKBUF_X1 G4319 (
	 );
   OAI221_X1 G4318 (
	 );
   INV_X1 G4317 (
	 );
   INV_X1 G4316 (
	 );
   AOI22_X1 G4315 (
	 );
   NOR2_X1 G4314 (
	 );
   CLKBUF_X1 G4313 (
	 );
   OAI211_X1 G4312 (
	 );
   INV_X1 G4311 (
	 );
   NAND4_X1 G4310 (
	 );
   NOR3_X1 G4309 (
	 );
   AND3_X1 G4308 (
	 );
   NOR2_X1 G4307 (
	 );
   OAI22_X1 G4306 (
	 );
   INV_X1 G4305 (
	 );
   INV_X1 G4304 (
	 );
   CLKBUF_X1 G4303 (
	 );
   CLKBUF_X1 G4302 (
	 );
   CLKBUF_X1 G4301 (
	 );
   CLKBUF_X1 G4300 (
	 );
   NOR2_X1 G4299 (
	 );
   AOI21_X1 G4298 (
	 );
   INV_X1 G4297 (
	 );
   MUX2_X1 G4296 (
	 );
   CLKBUF_X1 G4295 (
	 );
   CLKBUF_X1 G4294 (
	 );
   CLKBUF_X1 G4293 (
	 );
   CLKBUF_X1 G4292 (
	 );
   CLKBUF_X1 G4291 (
	 );
   OAI21_X1 G4290 (
	 );
   INV_X1 G4289 (
	 );
   NAND2_X1 G4288 (
	 );
   NAND2_X1 G4287 (
	 );
   OAI221_X1 G4286 (
	 );
   AOI22_X1 G4285 (
	 );
   CLKBUF_X1 G4284 (
	 );
   CLKBUF_X1 G4283 (
	 );
   CLKBUF_X1 G4282 (
	 );
   AND2_X1 G4281 (
	 );
   CLKBUF_X1 G4280 (
	 );
   AND2_X1 G4279 (
	 );
   NOR2_X1 G4278 (
	 );
   NAND2_X1 G4277 (
	 );
   AND4_X1 G4276 (
	 );
   NAND2_X1 G4275 (
	 );
   NAND2_X1 G4274 (
	 );
   NAND2_X1 G4273 (
	 );
   NAND2_X1 G4272 (
	 );
   AND4_X1 G4271 (
	 );
   NAND4_X1 G4270 (
	 );
   NAND4_X1 G4269 (
	 );
   NAND3_X1 G4268 (
	 );
   NAND3_X1 G4267 (
	 );
   CLKBUF_X1 G4266 (
	 );
   OAI21_X1 G4265 (
	 );
   INV_X1 G4264 (
	 );
   NAND2_X1 G4263 (
	 );
   MUX2_X1 G4262 (
	 );
   CLKBUF_X1 G4261 (
	 );
   CLKBUF_X1 G4260 (
	 );
   CLKBUF_X1 G4259 (
	 );
   CLKBUF_X1 G4258 (
	 );
   OAI21_X1 G4257 (
	 );
   INV_X1 G4256 (
	 );
   NAND2_X1 G4255 (
	 );
   CLKBUF_X1 G4254 (
	 );
   NAND2_X1 G4253 (
	 );
   AOI22_X1 G4252 (
	 );
   AOI22_X1 G4251 (
	 );
   NAND3_X1 G4250 (
	 );
   AOI22_X1 G4249 (
	 );
   AND3_X1 G4248 (
	 );
   NAND2_X1 G4247 (
	 );
   NAND2_X1 G4246 (
	 );
   NAND2_X1 G4245 (
	 );
   AND3_X1 G4244 (
	 );
   NAND4_X1 G4243 (
	 );
   NAND4_X1 G4242 (
	 );
   NAND4_X1 G4241 (
	 );
   OAI21_X1 G4240 (
	 );
   INV_X1 G4239 (
	 );
   NAND2_X1 G4238 (
	 );
   CLKBUF_X1 G4237 (
	 );
   CLKBUF_X1 G4236 (
	 );
   MUX2_X1 G4235 (
	 );
   OAI21_X1 G4234 (
	 );
   INV_X1 G4233 (
	 );
   NAND2_X1 G4232 (
	 );
   CLKBUF_X1 G4231 (
	 );
   CLKBUF_X1 G4230 (
	 );
   CLKBUF_X1 G4229 (
	 );
   CLKBUF_X1 G4228 (
	 );
   CLKBUF_X1 G4227 (
	 );
   OAI221_X1 G4226 (
	 );
   INV_X1 G4225 (
	 );
   AOI22_X1 G4224 (
	 );
   NAND3_X1 G4223 (
	 );
   AOI22_X1 G4222 (
	 );
   AND3_X1 G4221 (
	 );
   NAND2_X1 G4220 (
	 );
   NAND2_X1 G4219 (
	 );
   NAND2_X1 G4218 (
	 );
   AND3_X1 G4217 (
	 );
   NAND4_X1 G4216 (
	 );
   NAND4_X1 G4215 (
	 );
   NAND4_X1 G4214 (
	 );
   CLKBUF_X1 G4213 (
	 );
   CLKBUF_X1 G4212 (
	 );
   OAI21_X1 G4211 (
	 );
   INV_X1 G4210 (
	 );
   NAND2_X1 G4209 (
	 );
   CLKBUF_X1 G4208 (
	 );
   MUX2_X1 G4207 (
	 );
   MUX2_X1 G4206 (
	 );
   CLKBUF_X1 G4205 (
	 );
   NAND2_X1 G4204 (
	 );
   AOI22_X1 G4203 (
	 );
   AOI22_X1 G4202 (
	 );
   OAI21_X1 G4201 (
	 );
   INV_X1 G4200 (
	 );
   NAND2_X1 G4199 (
	 );
   NOR2_X1 G4198 (
	 );
   NAND2_X1 G4197 (
	 );
   AOI22_X1 G4196 (
	 );
   AOI22_X1 G4195 (
	 );
   CLKBUF_X1 G4194 (
	 );
   CLKBUF_X1 G4193 (
	 );
   CLKBUF_X1 G4192 (
	 );
   CLKBUF_X1 G4191 (
	 );
   CLKBUF_X1 G4190 (
	 );
   AOI21_X1 G4189 (
	 );
   INV_X1 G4188 (
	 );
   NOR2_X1 G4187 (
	 );
   CLKBUF_X1 G4186 (
	 );
   NAND3_X1 G4185 (
	 );
   AOI22_X1 G4184 (
	 );
   AND3_X1 G4183 (
	 );
   NAND2_X1 G4182 (
	 );
   NAND2_X1 G4181 (
	 );
   NAND2_X1 G4180 (
	 );
   AND3_X1 G4179 (
	 );
   NAND4_X1 G4178 (
	 );
   NAND4_X1 G4177 (
	 );
   NAND4_X1 G4176 (
	 );
   CLKBUF_X1 G4175 (
	 );
   NAND2_X1 G4174 (
	 );
   AOI22_X1 G4173 (
	 );
   AOI22_X1 G4172 (
	 );
   CLKBUF_X1 G4171 (
	 );
   CLKBUF_X1 G4170 (
	 );
   CLKBUF_X1 G4169 (
	 );
   MUX2_X1 G4168 (
	 );
   NAND2_X1 G4167 (
	 );
   AOI22_X1 G4166 (
	 );
   AOI22_X1 G4165 (
	 );
   OAI21_X1 G4164 (
	 );
   INV_X1 G4163 (
	 );
   NAND2_X1 G4162 (
	 );
   NAND2_X1 G4161 (
	 );
   NAND2_X1 G4160 (
	 );
   CLKBUF_X1 G4159 (
	 );
   MUX2_X1 G4158 (
	 );
   CLKBUF_X1 G4157 (
	 );
   CLKBUF_X1 G4156 (
	 );
   MUX2_X1 G4155 (
	 );
   CLKBUF_X1 G4154 (
	 );
   CLKBUF_X1 G4153 (
	 );
   CLKBUF_X1 G4152 (
	 );
   OAI21_X1 G4151 (
	 );
   INV_X1 G4150 (
	 );
   NAND2_X1 G4149 (
	 );
   CLKBUF_X1 G4148 (
	 );
   CLKBUF_X1 G4147 (
	 );
   OAI21_X1 G4146 (
	 );
   INV_X1 G4145 (
	 );
   NAND2_X1 G4144 (
	 );
   CLKBUF_X1 G4143 (
	 );
   AOI21_X1 G4142 (
	 );
   INV_X1 G4141 (
	 );
   NAND2_X1 G4140 (
	 );
   AND4_X1 G4139 (
	 );
   NAND2_X1 G4138 (
	 );
   NAND2_X1 G4137 (
	 );
   NAND2_X1 G4136 (
	 );
   NAND2_X1 G4135 (
	 );
   AND4_X1 G4134 (
	 );
   NAND4_X1 G4133 (
	 );
   NAND4_X1 G4132 (
	 );
   NAND3_X1 G4131 (
	 );
   NAND3_X1 G4130 (
	 );
   CLKBUF_X1 G4129 (
	 );
   NAND3_X1 G4128 (
	 );
   AOI22_X1 G4127 (
	 );
   AND3_X1 G4126 (
	 );
   NAND2_X1 G4125 (
	 );
   NAND2_X1 G4124 (
	 );
   NAND2_X1 G4123 (
	 );
   AND3_X1 G4122 (
	 );
   NAND4_X1 G4121 (
	 );
   NAND4_X1 G4120 (
	 );
   NAND4_X1 G4119 (
	 );
   CLKBUF_X1 G4118 (
	 );
   CLKBUF_X1 G4117 (
	 );
   CLKBUF_X1 G4116 (
	 );
   CLKBUF_X1 G4115 (
	 );
   CLKBUF_X1 G4114 (
	 );
   MUX2_X1 G4113 (
	 );
   CLKBUF_X1 G4112 (
	 );
   CLKBUF_X1 G4111 (
	 );
   NAND2_X1 G4110 (
	 );
   AND4_X1 G4109 (
	 );
   NAND2_X1 G4108 (
	 );
   NAND2_X1 G4107 (
	 );
   NAND4_X1 G4106 (
	 );
   NAND3_X1 G4105 (
	 );
   NAND3_X1 G4104 (
	 );
   NAND3_X1 G4103 (
	 );
   NAND2_X1 G4102 (
	 );
   NAND2_X1 G4101 (
	 );
   NAND4_X1 G4100 (
	 );
   NAND3_X1 G4099 (
	 );
   NAND3_X1 G4098 (
	 );
   NAND3_X1 G4097 (
	 );
   NAND2_X1 G4096 (
	 );
   NAND2_X1 G4095 (
	 );
   NAND4_X1 G4094 (
	 );
   NAND3_X1 G4093 (
	 );
   NAND3_X1 G4092 (
	 );
   NAND3_X1 G4091 (
	 );
   NAND2_X1 G4090 (
	 );
   AND4_X1 G4089 (
	 );
   NAND4_X1 G4088 (
	 );
   NAND4_X1 G4087 (
	 );
   NAND3_X1 G4086 (
	 );
   NAND3_X1 G4085 (
	 );
   CLKBUF_X1 G4084 (
	 );
   CLKBUF_X1 G4083 (
	 );
   AOI21_X1 G4082 (
	 );
   INV_X1 G4081 (
	 );
   NOR2_X1 G4080 (
	 );
   CLKBUF_X1 G4079 (
	 );
   CLKBUF_X1 G4078 (
	 );
   MUX2_X1 G4077 (
	 );
   NAND3_X1 G4076 (
	 );
   NAND4_X1 G4075 (
	 );
   NOR3_X1 G4074 (
	 );
   NAND3_X1 G4073 (
	 );
   NAND4_X1 G4072 (
	 );
   NAND3_X1 G4071 (
	 );
   NAND3_X1 G4070 (
	 );
   OAI22_X1 G4069 (
	 );
   INV_X1 G4068 (
	 );
   INV_X1 G4067 (
	 );
   AND4_X1 G4066 (
	 );
   NOR2_X1 G4065 (
	 );
   NOR2_X1 G4064 (
	 );
   NOR2_X1 G4063 (
	 );
   INV_X1 G4062 (
	 );
   CLKBUF_X1 G4061 (
	 );
   MUX2_X1 G4060 (
	 );
   CLKBUF_X1 G4059 (
	 );
   CLKBUF_X1 G4058 (
	 );
   CLKBUF_X1 G4057 (
	 );
   NAND4_X1 G4056 (
	 );
   NAND2_X1 G4055 (
	 );
   NAND2_X1 G4054 (
	 );
   NAND2_X1 G4053 (
	 );
   AOI22_X1 G4052 (
	 );
   AOI22_X1 G4051 (
	 );
   NAND2_X1 G4050 (
	 );
   NAND4_X1 G4049 (
	 );
   NAND3_X1 G4048 (
	 );
   NAND3_X1 G4047 (
	 );
   NAND3_X1 G4046 (
	 );
   NAND2_X1 G4045 (
	 );
   AOI22_X1 G4044 (
	 );
   CLKBUF_X1 G4043 (
	 );
   AND2_X1 G4042 (
	 );
   MUX2_X1 G4041 (
	 );
   CLKBUF_X1 G4040 (
	 );
   CLKBUF_X1 G4039 (
	 );
   NAND4_X1 G4038 (
	 );
   AOI22_X1 G4037 (
	 );
   NAND2_X1 G4036 (
	 );
   NAND2_X1 G4035 (
	 );
   NAND2_X1 G4034 (
	 );
   CLKBUF_X1 G4033 (
	 );
   OAI221_X1 G4032 (
	 );
   AOI22_X1 G4031 (
	 );
   CLKBUF_X1 G4030 (
	 );
   CLKBUF_X1 G4029 (
	 );
   CLKBUF_X1 G4028 (
	 );
   NOR2_X1 G4027 (
	 );
   XNOR2_X1 G4026 (
	 );
   NAND4_X1 G4025 (
	 );
   NAND3_X1 G4024 (
	 );
   NAND2_X1 G4023 (
	 );
   NAND2_X1 G4022 (
	 );
   OAI21_X1 G4021 (
	 );
   OAI21_X1 G4020 (
	 );
   INV_X1 G4019 (
	 );
   NAND2_X1 G4018 (
	 );
   NAND2_X1 G4017 (
	 );
   AND4_X1 G4016 (
	 );
   NAND2_X1 G4015 (
	 );
   NAND2_X1 G4014 (
	 );
   NAND2_X1 G4013 (
	 );
   NAND2_X1 G4012 (
	 );
   NAND4_X1 G4011 (
	 );
   NAND3_X1 G4010 (
	 );
   NAND3_X1 G4009 (
	 );
   NAND3_X1 G4008 (
	 );
   NAND2_X1 G4007 (
	 );
   AND4_X1 G4006 (
	 );
   NAND4_X1 G4005 (
	 );
   NAND4_X1 G4004 (
	 );
   NAND3_X1 G4003 (
	 );
   NAND3_X1 G4002 (
	 );
   OAI221_X1 G4001 (
	 );
   INV_X1 G4000 (
	 );
   AOI22_X1 G3999 (
	 );
   CLKBUF_X1 G3998 (
	 );
   AOI21_X1 G3997 (
	 );
   NAND3_X1 G3996 (
	 );
   NOR2_X1 G3995 (
	 );
   CLKBUF_X1 G3994 (
	 );
   NOR2_X1 G3993 (
	 );
   NAND2_X1 G3992 (
	 );
   NAND2_X1 G3991 (
	 );
   AOI22_X1 G3990 (
	 );
   CLKBUF_X1 G3989 (
	 );
   CLKBUF_X1 G3988 (
	 );
   MUX2_X1 G3987 (
	 );
   CLKBUF_X1 G3986 (
	 );
   CLKBUF_X1 G3985 (
	 );
   MUX2_X1 G3984 (
	 );
   NAND2_X1 G3983 (
	 );
   NAND2_X1 G3982 (
	 );
   AOI22_X1 G3981 (
	 );
   AND2_X1 G3980 (
	 );
   CLKBUF_X1 G3979 (
	 );
   AOI21_X1 G3978 (
	 );
   INV_X1 G3977 (
	 );
   NAND3_X1 G3976 (
	 );
   AOI21_X1 G3975 (
	 );
   AOI21_X1 G3974 (
	 );
   OAI21_X1 G3973 (
	 );
   INV_X1 G3972 (
	 );
   NOR2_X1 G3971 (
	 );
   CLKBUF_X1 G3970 (
	 );
   CLKBUF_X1 G3969 (
	 );
   CLKBUF_X1 G3968 (
	 );
   CLKBUF_X1 G3967 (
	 );
   CLKBUF_X1 G3966 (
	 );
   CLKBUF_X1 G3965 (
	 );
   CLKBUF_X1 G3964 (
	 );
   OAI221_X1 G3963 (
	 );
   INV_X1 G3962 (
	 );
   INV_X1 G3961 (
	 );
   AOI22_X1 G3960 (
	 );
   CLKBUF_X1 G3959 (
	 );
   CLKBUF_X1 G3958 (
	 );
   CLKBUF_X1 G3957 (
	 );
   CLKBUF_X1 G3956 (
	 );
   CLKBUF_X1 G3955 (
	 );
   CLKBUF_X1 G3954 (
	 );
   CLKBUF_X1 G3953 (
	 );
   CLKBUF_X1 G3952 (
	 );
   OAI21_X1 G3951 (
	 );
   INV_X1 G3950 (
	 );
   NAND2_X1 G3949 (
	 );
   NOR3_X1 G3948 (
	 );
   AOI21_X1 G3947 (
	 );
   CLKBUF_X1 G3946 (
	 );
   CLKBUF_X1 G3945 (
	 );
   OAI221_X1 G3944 (
	 );
   INV_X1 G3943 (
	 );
   AOI22_X1 G3942 (
	 );
   NOR2_X1 G3941 (
	 );
   CLKBUF_X1 G3940 (
	 );
   CLKBUF_X1 G3939 (
	 );
   CLKBUF_X1 G3938 (
	 );
   OAI21_X1 G3937 (
	 );
   INV_X1 G3936 (
	 );
   NAND2_X1 G3935 (
	 );
   CLKBUF_X1 G3934 (
	 );
   CLKBUF_X1 G3933 (
	 );
   CLKBUF_X1 G3932 (
	 );
   NAND3_X1 G3931 (
	 );
   AOI22_X1 G3930 (
	 );
   AND3_X1 G3929 (
	 );
   NAND2_X1 G3928 (
	 );
   NAND2_X1 G3927 (
	 );
   NAND2_X1 G3926 (
	 );
   NAND4_X1 G3925 (
	 );
   NAND3_X1 G3924 (
	 );
   NAND3_X1 G3923 (
	 );
   NAND3_X1 G3922 (
	 );
   NAND2_X1 G3921 (
	 );
   AND3_X1 G3920 (
	 );
   NAND4_X1 G3919 (
	 );
   NAND4_X1 G3918 (
	 );
   NAND4_X1 G3917 (
	 );
   CLKBUF_X1 G3916 (
	 );
   CLKBUF_X1 G3915 (
	 );
   MUX2_X1 G3914 (
	 );
   AOI21_X1 G3913 (
	 );
   OAI21_X1 G3912 (
	 );
   NOR3_X1 G3911 (
	 );
   INV_X1 G3910 (
	 );
   CLKBUF_X1 G3909 (
	 );
   OAI21_X1 G3908 (
	 );
   INV_X1 G3907 (
	 );
   NAND2_X1 G3906 (
	 );
   CLKBUF_X1 G3905 (
	 );
   CLKBUF_X1 G3904 (
	 );
   CLKBUF_X1 G3903 (
	 );
   OAI21_X1 G3902 (
	 );
   NAND2_X1 G3901 (
	 );
   CLKBUF_X1 G3900 (
	 );
   NAND3_X1 G3899 (
	 );
   AND3_X1 G3898 (
	 );
   NAND2_X1 G3897 (
	 );
   NAND2_X1 G3896 (
	 );
   NAND4_X1 G3895 (
	 );
   NAND3_X1 G3894 (
	 );
   NAND3_X1 G3893 (
	 );
   NAND3_X1 G3892 (
	 );
   NAND2_X1 G3891 (
	 );
   NAND2_X1 G3890 (
	 );
   AOI22_X1 G3889 (
	 );
   AND3_X1 G3888 (
	 );
   NAND4_X1 G3887 (
	 );
   NAND4_X1 G3886 (
	 );
   NAND4_X1 G3885 (
	 );
   CLKBUF_X1 G3884 (
	 );
   CLKBUF_X1 G3883 (
	 );
   MUX2_X1 G3882 (
	 );
   CLKBUF_X1 G3881 (
	 );
   CLKBUF_X1 G3880 (
	 );
   OAI21_X1 G3879 (
	 );
   NAND2_X1 G3878 (
	 );
   OAI21_X1 G3877 (
	 );
   NOR2_X1 G3876 (
	 );
   NOR2_X1 G3875 (
	 );
   CLKBUF_X1 G3874 (
	 );
   NOR2_X1 G3873 (
	 );
   CLKBUF_X1 G3872 (
	 );
   NOR3_X1 G3871 (
	 );
   NOR2_X1 G3870 (
	 );
   AND2_X1 G3869 (
	 );
   AND2_X1 G3868 (
	 );
   NOR2_X1 G3867 (
	 );
   NAND3_X1 G3866 (
	 );
   OR2_X1 G3865 (
	 );
   NOR3_X1 G3864 (
	 );
   NAND3_X1 G3863 (
	 );
   NAND4_X1 G3862 (
	 );
   NAND3_X1 G3861 (
	 );
   NAND3_X1 G3860 (
	 );
   OAI22_X1 G3859 (
	 );
   INV_X1 G3858 (
	 );
   INV_X1 G3857 (
	 );
   AND4_X1 G3856 (
	 );
   NOR2_X1 G3855 (
	 );
   NOR2_X1 G3854 (
	 );
   NOR2_X1 G3853 (
	 );
   INV_X1 G3852 (
	 );
   CLKBUF_X1 G3851 (
	 );
   OAI221_X1 G3850 (
	 );
   AOI22_X1 G3849 (
	 );
   CLKBUF_X1 G3848 (
	 );
   OAI221_X1 G3847 (
	 );
   INV_X1 G3846 (
	 );
   AOI22_X1 G3845 (
	 );
   OAI21_X1 G3844 (
	 );
   INV_X1 G3843 (
	 );
   NAND2_X1 G3842 (
	 );
   CLKBUF_X1 G3841 (
	 );
   CLKBUF_X1 G3840 (
	 );
   CLKBUF_X1 G3839 (
	 );
   OAI221_X1 G3838 (
	 );
   INV_X1 G3837 (
	 );
   AOI22_X1 G3836 (
	 );
   OAI221_X1 G3835 (
	 );
   AOI22_X1 G3834 (
	 );
   CLKBUF_X1 G3833 (
	 );
   CLKBUF_X1 G3832 (
	 );
   NAND2_X1 G3831 (
	 );
   OAI221_X1 G3830 (
	 );
   INV_X1 G3829 (
	 );
   INV_X1 G3828 (
	 );
   AOI22_X1 G3827 (
	 );
   BUF_X4 G3826 (
	 );
   BUF_X4 G3825 (
	 );
   NOR2_X1 G3824 (
	 );
   NAND3_X1 G3823 (
	 );
   AOI22_X1 G3822 (
	 );
   AND3_X1 G3821 (
	 );
   NAND2_X1 G3820 (
	 );
   NAND2_X1 G3819 (
	 );
   NAND2_X1 G3818 (
	 );
   NAND4_X1 G3817 (
	 );
   NAND3_X1 G3816 (
	 );
   NAND3_X1 G3815 (
	 );
   NAND3_X1 G3814 (
	 );
   NAND2_X1 G3813 (
	 );
   AND3_X1 G3812 (
	 );
   NAND4_X1 G3811 (
	 );
   NAND4_X1 G3810 (
	 );
   NAND4_X1 G3809 (
	 );
   CLKBUF_X1 G3808 (
	 );
   OAI21_X1 G3807 (
	 );
   INV_X1 G3806 (
	 );
   NAND2_X1 G3805 (
	 );
   CLKBUF_X1 G3804 (
	 );
   MUX2_X1 G3803 (
	 );
   CLKBUF_X1 G3802 (
	 );
   NAND4_X1 G3801 (
	 );
   NAND2_X1 G3800 (
	 );
   NAND2_X1 G3799 (
	 );
   NAND2_X1 G3798 (
	 );
   AOI22_X1 G3797 (
	 );
   NAND2_X1 G3796 (
	 );
   AOI22_X1 G3795 (
	 );
   AOI22_X1 G3794 (
	 );
   OAI21_X1 G3793 (
	 );
   INV_X1 G3792 (
	 );
   NAND2_X1 G3791 (
	 );
   CLKBUF_X1 G3790 (
	 );
   CLKBUF_X1 G3789 (
	 );
   NAND4_X1 G3788 (
	 );
   AOI22_X1 G3787 (
	 );
   NAND2_X1 G3786 (
	 );
   NAND2_X1 G3785 (
	 );
   NAND2_X1 G3784 (
	 );
   AND2_X1 G3783 (
	 );
   CLKBUF_X1 G3782 (
	 );
   CLKBUF_X1 G3781 (
	 );
   AND2_X1 G3780 (
	 );
   CLKBUF_X1 G3779 (
	 );
   CLKBUF_X1 G3778 (
	 );
   NOR3_X1 G3777 (
	 );
   AOI21_X1 G3776 (
	 );
   NOR3_X1 G3775 (
	 );
   CLKBUF_X1 G3774 (
	 );
   CLKBUF_X1 G3773 (
	 );
   CLKBUF_X1 G3772 (
	 );
   AOI21_X1 G3771 (
	 );
   NAND3_X1 G3770 (
	 );
   AOI22_X1 G3769 (
	 );
   AND3_X1 G3768 (
	 );
   NAND2_X1 G3767 (
	 );
   NAND2_X1 G3766 (
	 );
   NAND4_X1 G3765 (
	 );
   NAND3_X1 G3764 (
	 );
   NAND3_X1 G3763 (
	 );
   NAND3_X1 G3762 (
	 );
   NAND2_X1 G3761 (
	 );
   NAND2_X1 G3760 (
	 );
   AND3_X1 G3759 (
	 );
   NAND4_X1 G3758 (
	 );
   NAND4_X1 G3757 (
	 );
   NAND4_X1 G3756 (
	 );
   CLKBUF_X1 G3755 (
	 );
   AND2_X1 G3754 (
	 );
   CLKBUF_X1 G3753 (
	 );
   CLKBUF_X1 G3752 (
	 );
   CLKBUF_X1 G3751 (
	 );
   OAI21_X1 G3750 (
	 );
   INV_X1 G3749 (
	 );
   NAND2_X1 G3748 (
	 );
   NOR2_X1 G3747 (
	 );
   NAND4_X1 G3746 (
	 );
   NAND4_X1 G3745 (
	 );
   NAND2_X1 G3744 (
	 );
   AOI22_X1 G3743 (
	 );
   AOI22_X1 G3742 (
	 );
   CLKBUF_X1 G3741 (
	 );
   AOI21_X1 G3740 (
	 );
   OAI21_X1 G3739 (
	 );
   AND3_X1 G3738 (
	 );
   CLKBUF_X1 G3737 (
	 );
   CLKBUF_X1 G3736 (
	 );
   OAI21_X1 G3735 (
	 );
   INV_X1 G3734 (
	 );
   NAND2_X1 G3733 (
	 );
   CLKBUF_X1 G3732 (
	 );
   NAND3_X1 G3731 (
	 );
   AOI22_X1 G3730 (
	 );
   AND3_X1 G3729 (
	 );
   NAND2_X1 G3728 (
	 );
   NAND2_X1 G3727 (
	 );
   NAND2_X1 G3726 (
	 );
   AND3_X1 G3725 (
	 );
   NAND4_X1 G3724 (
	 );
   NAND4_X1 G3723 (
	 );
   NAND4_X1 G3722 (
	 );
   CLKBUF_X1 G3721 (
	 );
   CLKBUF_X1 G3720 (
	 );
   NAND2_X1 G3719 (
	 );
   AOI22_X1 G3718 (
	 );
   AOI22_X1 G3717 (
	 );
   CLKBUF_X1 G3716 (
	 );
   NAND3_X1 G3715 (
	 );
   AND3_X1 G3714 (
	 );
   NAND2_X1 G3713 (
	 );
   NAND2_X1 G3712 (
	 );
   NAND2_X1 G3711 (
	 );
   AOI22_X1 G3710 (
	 );
   AND3_X1 G3709 (
	 );
   NAND4_X1 G3708 (
	 );
   NAND4_X1 G3707 (
	 );
   NAND4_X1 G3706 (
	 );
   MUX2_X1 G3705 (
	 );
   CLKBUF_X1 G3704 (
	 );
   CLKBUF_X1 G3703 (
	 );
   CLKBUF_X1 G3702 (
	 );
   CLKBUF_X1 G3701 (
	 );
   CLKBUF_X1 G3700 (
	 );
   NAND2_X1 G3699 (
	 );
   NAND2_X1 G3698 (
	 );
   AOI22_X1 G3697 (
	 );
   OAI21_X1 G3696 (
	 );
   INV_X1 G3695 (
	 );
   NAND2_X1 G3694 (
	 );
   OAI21_X1 G3693 (
	 );
   NOR2_X1 G3692 (
	 );
   NOR2_X1 G3691 (
	 );
   OAI221_X1 G3690 (
	 );
   NAND2_X1 G3689 (
	 );
   OAI21_X1 G3688 (
	 );
   OAI21_X1 G3687 (
	 );
   CLKBUF_X1 G3686 (
	 );
   OAI21_X1 G3685 (
	 );
   INV_X1 G3684 (
	 );
   NAND2_X1 G3683 (
	 );
   CLKBUF_X1 G3682 (
	 );
   CLKBUF_X1 G3681 (
	 );
   MUX2_X1 G3680 (
	 );
   CLKBUF_X1 G3679 (
	 );
   CLKBUF_X1 G3678 (
	 );
   CLKBUF_X1 G3677 (
	 );
   CLKBUF_X1 G3676 (
	 );
   MUX2_X1 G3675 (
	 );
   CLKBUF_X1 G3674 (
	 );
   CLKBUF_X1 G3673 (
	 );
   MUX2_X1 G3672 (
	 );
   CLKBUF_X1 G3671 (
	 );
   CLKBUF_X1 G3670 (
	 );
   CLKBUF_X1 G3669 (
	 );
   CLKBUF_X1 G3668 (
	 );
   CLKBUF_X1 G3667 (
	 );
   OAI21_X1 G3666 (
	 );
   INV_X1 G3665 (
	 );
   NAND2_X1 G3664 (
	 );
   CLKBUF_X1 G3663 (
	 );
   MUX2_X1 G3662 (
	 );
   XNOR2_X1 G3661 (
	 );
   NAND2_X1 G3660 (
	 );
   XNOR2_X1 G3659 (
	 );
   CLKBUF_X1 G3658 (
	 );
   CLKBUF_X1 G3657 (
	 );
   CLKBUF_X1 G3656 (
	 );
   AND2_X1 G3655 (
	 );
   CLKBUF_X1 G3654 (
	 );
   CLKBUF_X1 G3653 (
	 );
   NOR2_X1 G3652 (
	 );
   AOI21_X1 G3651 (
	 );
   INV_X1 G3650 (
	 );
   INV_X1 G3649 (
	 );
   NAND2_X1 G3648 (
	 );
   AOI22_X1 G3647 (
	 );
   AOI22_X1 G3646 (
	 );
   CLKBUF_X1 G3645 (
	 );
   CLKBUF_X1 G3644 (
	 );
   CLKBUF_X1 G3643 (
	 );
   OAI221_X1 G3642 (
	 );
   AOI22_X1 G3641 (
	 );
   CLKBUF_X1 G3640 (
	 );
   NAND2_X1 G3639 (
	 );
   AOI22_X1 G3638 (
	 );
   AOI22_X1 G3637 (
	 );
   AND2_X1 G3636 (
	 );
   MUX2_X1 G3635 (
	 );
   BUF_X8 G3634 (
	 );
   CLKBUF_X1 G3633 (
	 );
   CLKBUF_X1 G3632 (
	 );
   CLKBUF_X1 G3631 (
	 );
   NOR2_X1 G3630 (
	 );
   INV_X1 G3629 (
	 );
   CLKBUF_X1 G3628 (
	 );
   CLKBUF_X1 G3627 (
	 );
   CLKBUF_X1 G3626 (
	 );
   NAND3_X1 G3625 (
	 );
   AOI22_X1 G3624 (
	 );
   AND3_X1 G3623 (
	 );
   NAND2_X1 G3622 (
	 );
   NAND2_X1 G3621 (
	 );
   NAND2_X1 G3620 (
	 );
   AND3_X1 G3619 (
	 );
   NAND4_X1 G3618 (
	 );
   NAND4_X1 G3617 (
	 );
   NAND4_X1 G3616 (
	 );
   CLKBUF_X1 G3615 (
	 );
   CLKBUF_X1 G3614 (
	 );
   CLKBUF_X1 G3613 (
	 );
   CLKBUF_X1 G3612 (
	 );
   OAI22_X1 G3611 (
	 );
   OAI21_X1 G3610 (
	 );
   XNOR2_X1 G3609 (
	 );
   OAI21_X1 G3608 (
	 );
   XNOR2_X1 G3607 (
	 );
   INV_X1 G3606 (
	 );
   AOI22_X1 G3605 (
	 );
   CLKBUF_X1 G3604 (
	 );
   MUX2_X1 G3603 (
	 );
   CLKBUF_X1 G3602 (
	 );
   CLKBUF_X1 G3601 (
	 );
   CLKBUF_X1 G3600 (
	 );
   MUX2_X1 G3599 (
	 );
   CLKBUF_X1 G3598 (
	 );
   CLKBUF_X1 G3597 (
	 );
   INV_X1 G3596 (
	 );
   NAND2_X1 G3595 (
	 );
   CLKBUF_X1 G3594 (
	 );
   OAI221_X1 G3593 (
	 );
   AOI22_X1 G3592 (
	 );
   CLKBUF_X1 G3591 (
	 );
   AND2_X1 G3590 (
	 );
   CLKBUF_X1 G3589 (
	 );
   CLKBUF_X1 G3588 (
	 );
   CLKBUF_X1 G3587 (
	 );
   MUX2_X1 G3586 (
	 );
   AOI21_X1 G3585 (
	 );
   OAI21_X1 G3584 (
	 );
   CLKBUF_X1 G3583 (
	 );
   AND3_X1 G3582 (
	 );
   CLKBUF_X1 G3581 (
	 );
   CLKBUF_X1 G3580 (
	 );
   CLKBUF_X1 G3579 (
	 );
   MUX2_X1 G3578 (
	 );
   AND2_X1 G3577 (
	 );
   AOI21_X1 G3576 (
	 );
   INV_X1 G3575 (
	 );
   NAND3_X1 G3574 (
	 );
   AOI22_X1 G3573 (
	 );
   AND3_X1 G3572 (
	 );
   NAND2_X1 G3571 (
	 );
   NAND2_X1 G3570 (
	 );
   NAND4_X1 G3569 (
	 );
   NAND3_X1 G3568 (
	 );
   NAND3_X1 G3567 (
	 );
   NAND3_X1 G3566 (
	 );
   NAND2_X1 G3565 (
	 );
   NAND2_X1 G3564 (
	 );
   AND3_X1 G3563 (
	 );
   NAND4_X1 G3562 (
	 );
   NAND4_X1 G3561 (
	 );
   NAND4_X1 G3560 (
	 );
   CLKBUF_X1 G3559 (
	 );
   CLKBUF_X1 G3558 (
	 );
   CLKBUF_X1 G3557 (
	 );
   CLKBUF_X1 G3556 (
	 );
   OAI21_X1 G3555 (
	 );
   INV_X1 G3554 (
	 );
   NAND2_X1 G3553 (
	 );
   NAND3_X1 G3552 (
	 );
   AOI22_X1 G3551 (
	 );
   AND3_X1 G3550 (
	 );
   NAND2_X1 G3549 (
	 );
   NAND2_X1 G3548 (
	 );
   NAND2_X1 G3547 (
	 );
   AND3_X1 G3546 (
	 );
   NAND4_X1 G3545 (
	 );
   NAND4_X1 G3544 (
	 );
   NAND4_X1 G3543 (
	 );
   AND2_X1 G3542 (
	 );
   CLKBUF_X1 G3541 (
	 );
   CLKBUF_X1 G3540 (
	 );
   MUX2_X1 G3539 (
	 );
   CLKBUF_X1 G3538 (
	 );
   OAI21_X1 G3537 (
	 );
   INV_X1 G3536 (
	 );
   NAND2_X1 G3535 (
	 );
   AOI21_X1 G3534 (
	 );
   INV_X1 G3533 (
	 );
   NOR2_X1 G3532 (
	 );
   AND2_X1 G3531 (
	 );
   CLKBUF_X1 G3530 (
	 );
   CLKBUF_X1 G3529 (
	 );
   NOR2_X1 G3528 (
	 );
   CLKBUF_X1 G3527 (
	 );
   MUX2_X1 G3526 (
	 );
   CLKBUF_X1 G3525 (
	 );
   AOI21_X1 G3524 (
	 );
   NAND3_X1 G3523 (
	 );
   INV_X1 G3522 (
	 );
   AND2_X1 G3521 (
	 );
   INV_X1 G3520 (
	 );
   AOI211_X1 G3519 (
	 );
   AOI21_X1 G3518 (
	 );
   OAI21_X1 G3517 (
	 );
   INV_X1 G3516 (
	 );
   NOR2_X1 G3515 (
	 );
   INV_X1 G3514 (
	 );
   OAI211_X1 G3513 (
	 );
   INV_X1 G3512 (
	 );
   NAND2_X1 G3511 (
	 );
   AOI21_X1 G3510 (
	 );
   OAI22_X1 G3509 (
	 );
   INV_X1 G3508 (
	 );
   INV_X1 G3507 (
	 );
   CLKBUF_X1 G3506 (
	 );
   NAND4_X1 G3505 (
	 );
   NAND4_X1 G3504 (
	 );
   OR2_X1 G3503 (
	 );
   NAND4_X1 G3502 (
	 );
   NOR2_X1 G3501 (
	 );
   AND2_X1 G3500 (
	 );
   NAND4_X1 G3499 (
	 );
   NAND4_X1 G3498 (
	 );
   NAND3_X1 G3497 (
	 );
   NAND3_X1 G3496 (
	 );
   NAND4_X1 G3495 (
	 );
   CLKBUF_X1 G3494 (
	 );
   OAI21_X1 G3493 (
	 );
   INV_X1 G3492 (
	 );
   NAND2_X1 G3491 (
	 );
   CLKBUF_X1 G3490 (
	 );
   CLKBUF_X1 G3489 (
	 );
   MUX2_X1 G3488 (
	 );
   OAI21_X1 G3487 (
	 );
   INV_X1 G3486 (
	 );
   NAND2_X1 G3485 (
	 );
   CLKBUF_X1 G3484 (
	 );
   CLKBUF_X1 G3483 (
	 );
   MUX2_X1 G3482 (
	 );
   AND2_X1 G3481 (
	 );
   CLKBUF_X1 G3480 (
	 );
   NOR2_X1 G3479 (
	 );
   CLKBUF_X1 G3478 (
	 );
   MUX2_X1 G3477 (
	 );
   CLKBUF_X1 G3476 (
	 );
   MUX2_X1 G3475 (
	 );
   CLKBUF_X1 G3474 (
	 );
   CLKBUF_X1 G3473 (
	 );
   CLKBUF_X1 G3472 (
	 );
   MUX2_X1 G3471 (
	 );
   CLKBUF_X1 G3470 (
	 );
   OAI21_X1 G3469 (
	 );
   INV_X1 G3468 (
	 );
   NAND2_X1 G3467 (
	 );
   CLKBUF_X1 G3466 (
	 );
   MUX2_X1 G3465 (
	 );
   AOI21_X1 G3464 (
	 );
   INV_X1 G3463 (
	 );
   NOR2_X1 G3462 (
	 );
   CLKBUF_X1 G3461 (
	 );
   OAI221_X1 G3460 (
	 );
   INV_X1 G3459 (
	 );
   AOI22_X1 G3458 (
	 );
   CLKBUF_X1 G3457 (
	 );
   NAND3_X1 G3456 (
	 );
   AOI22_X1 G3455 (
	 );
   AND3_X1 G3454 (
	 );
   NAND2_X1 G3453 (
	 );
   NAND2_X1 G3452 (
	 );
   NAND4_X1 G3451 (
	 );
   NAND3_X1 G3450 (
	 );
   NAND3_X1 G3449 (
	 );
   NAND3_X1 G3448 (
	 );
   NAND2_X1 G3447 (
	 );
   NAND2_X1 G3446 (
	 );
   AND3_X1 G3445 (
	 );
   NAND4_X1 G3444 (
	 );
   NAND4_X1 G3443 (
	 );
   NAND4_X1 G3442 (
	 );
   CLKBUF_X1 G3441 (
	 );
   CLKBUF_X1 G3440 (
	 );
   CLKBUF_X1 G3439 (
	 );
   MUX2_X1 G3438 (
	 );
   CLKBUF_X1 G3437 (
	 );
   CLKBUF_X1 G3436 (
	 );
   CLKBUF_X1 G3435 (
	 );
   AOI21_X1 G3434 (
	 );
   INV_X1 G3433 (
	 );
   NOR2_X1 G3432 (
	 );
   CLKBUF_X1 G3431 (
	 );
   OAI21_X1 G3430 (
	 );
   NAND2_X1 G3429 (
	 );
   NAND3_X1 G3428 (
	 );
   OAI21_X1 G3427 (
	 );
   CLKBUF_X1 G3426 (
	 );
   CLKBUF_X1 G3425 (
	 );
   MUX2_X1 G3424 (
	 );
   CLKBUF_X1 G3423 (
	 );
   AOI21_X1 G3422 (
	 );
   NAND2_X1 G3421 (
	 );
   OR2_X1 G3420 (
	 );
   AOI21_X1 G3419 (
	 );
   NAND3_X1 G3418 (
	 );
   INV_X1 G3417 (
	 );
   CLKBUF_X1 G3416 (
	 );
   OAI21_X1 G3415 (
	 );
   INV_X1 G3414 (
	 );
   NAND2_X1 G3413 (
	 );
   CLKBUF_X1 G3412 (
	 );
   CLKBUF_X1 G3411 (
	 );
   MUX2_X1 G3410 (
	 );
   CLKBUF_X1 G3409 (
	 );
   AND2_X1 G3408 (
	 );
   AOI21_X1 G3407 (
	 );
   INV_X1 G3406 (
	 );
   INV_X1 G3405 (
	 );
   OAI21_X1 G3404 (
	 );
   INV_X1 G3403 (
	 );
   NAND2_X1 G3402 (
	 );
   OAI21_X1 G3401 (
	 );
   INV_X1 G3400 (
	 );
   AOI22_X1 G3399 (
	 );
   CLKBUF_X1 G3398 (
	 );
   OAI21_X1 G3397 (
	 );
   INV_X1 G3396 (
	 );
   NAND2_X1 G3395 (
	 );
   CLKBUF_X1 G3394 (
	 );
   MUX2_X1 G3393 (
	 );
   OAI21_X1 G3392 (
	 );
   NAND2_X1 G3391 (
	 );
   CLKBUF_X1 G3390 (
	 );
   CLKBUF_X1 G3389 (
	 );
   CLKBUF_X1 G3388 (
	 );
   CLKBUF_X1 G3387 (
	 );
   AOI21_X1 G3386 (
	 );
   INV_X1 G3385 (
	 );
   NOR2_X1 G3384 (
	 );
   MUX2_X1 G3383 (
	 );
   OAI21_X1 G3382 (
	 );
   INV_X1 G3381 (
	 );
   AOI22_X1 G3380 (
	 );
   CLKBUF_X1 G3379 (
	 );
   CLKBUF_X1 G3378 (
	 );
   NAND2_X1 G3377 (
	 );
   AND4_X1 G3376 (
	 );
   NAND2_X1 G3375 (
	 );
   NAND2_X1 G3374 (
	 );
   NAND2_X1 G3373 (
	 );
   NAND2_X1 G3372 (
	 );
   AND4_X1 G3371 (
	 );
   NAND4_X1 G3370 (
	 );
   NAND4_X1 G3369 (
	 );
   NAND3_X1 G3368 (
	 );
   NAND3_X1 G3367 (
	 );
   OAI221_X1 G3366 (
	 );
   XNOR2_X1 G3365 (
	 );
   NAND3_X1 G3364 (
	 );
   NAND2_X1 G3363 (
	 );
   NAND4_X1 G3362 (
	 );
   OAI21_X1 G3361 (
	 );
   INV_X1 G3360 (
	 );
   NAND2_X1 G3359 (
	 );
   CLKBUF_X1 G3358 (
	 );
   OAI21_X1 G3357 (
	 );
   INV_X1 G3356 (
	 );
   INV_X1 G3355 (
	 );
   NAND2_X1 G3354 (
	 );
   CLKBUF_X1 G3353 (
	 );
   CLKBUF_X1 G3352 (
	 );
   CLKBUF_X1 G3351 (
	 );
   CLKBUF_X1 G3350 (
	 );
   CLKBUF_X1 G3349 (
	 );
   CLKBUF_X1 G3348 (
	 );
   OAI21_X1 G3347 (
	 );
   INV_X1 G3346 (
	 );
   NAND2_X1 G3345 (
	 );
   MUX2_X1 G3344 (
	 );
   CLKBUF_X1 G3343 (
	 );
   CLKBUF_X1 G3342 (
	 );
   CLKBUF_X1 G3341 (
	 );
   CLKBUF_X1 G3340 (
	 );
   AOI21_X1 G3339 (
	 );
   INV_X1 G3338 (
	 );
   NOR2_X1 G3337 (
	 );
   CLKBUF_X1 G3336 (
	 );
   NAND2_X1 G3335 (
	 );
   AOI22_X1 G3334 (
	 );
   AOI22_X1 G3333 (
	 );
   AOI211_X1 G3332 (
	 );
   CLKBUF_X1 G3331 (
	 );
   CLKBUF_X1 G3330 (
	 );
   NOR2_X1 G3329 (
	 );
   INV_X1 G3328 (
	 );
   NOR3_X1 G3327 (
	 );
   INV_X1 G3326 (
	 );
   AOI21_X1 G3325 (
	 );
   AND3_X1 G3324 (
	 );
   NOR2_X1 G3323 (
	 );
   INV_X1 G3322 (
	 );
   NAND2_X1 G3321 (
	 );
   OAI221_X1 G3320 (
	 );
   AOI22_X1 G3319 (
	 );
   NAND4_X1 G3318 (
	 );
   NAND4_X1 G3317 (
	 );
   OR2_X1 G3316 (
	 );
   OR2_X1 G3315 (
	 );
   NOR2_X1 G3314 (
	 );
   AND2_X1 G3313 (
	 );
   NAND4_X1 G3312 (
	 );
   NAND4_X1 G3311 (
	 );
   NAND3_X1 G3310 (
	 );
   NAND3_X1 G3309 (
	 );
   NAND4_X1 G3308 (
	 );
   CLKBUF_X1 G3307 (
	 );
   OAI21_X1 G3306 (
	 );
   INV_X1 G3305 (
	 );
   NAND2_X1 G3304 (
	 );
   CLKBUF_X1 G3303 (
	 );
   AOI21_X1 G3302 (
	 );
   NAND3_X1 G3301 (
	 );
   INV_X1 G3300 (
	 );
   OAI21_X1 G3299 (
	 );
   INV_X1 G3298 (
	 );
   NAND2_X1 G3297 (
	 );
   OAI21_X1 G3296 (
	 );
   NAND2_X1 G3295 (
	 );
   CLKBUF_X1 G3294 (
	 );
   CLKBUF_X1 G3293 (
	 );
   OAI21_X1 G3292 (
	 );
   NAND2_X1 G3291 (
	 );
   NOR2_X1 G3290 (
	 );
   CLKBUF_X1 G3289 (
	 );
   NOR2_X1 G3288 (
	 );
   CLKBUF_X1 G3287 (
	 );
   MUX2_X1 G3286 (
	 );
   CLKBUF_X1 G3285 (
	 );
   CLKBUF_X1 G3284 (
	 );
   NOR2_X1 G3283 (
	 );
   CLKBUF_X1 G3282 (
	 );
   AOI21_X1 G3281 (
	 );
   OAI21_X1 G3280 (
	 );
   NOR3_X1 G3279 (
	 );
   INV_X1 G3278 (
	 );
   AOI21_X1 G3277 (
	 );
   INV_X1 G3276 (
	 );
   INV_X1 G3275 (
	 );
   CLKBUF_X1 G3274 (
	 );
   CLKBUF_X1 G3273 (
	 );
   CLKBUF_X1 G3272 (
	 );
   CLKBUF_X1 G3271 (
	 );
   NAND3_X1 G3270 (
	 );
   AND3_X1 G3269 (
	 );
   NAND2_X1 G3268 (
	 );
   NAND4_X1 G3267 (
	 );
   NAND2_X1 G3266 (
	 );
   INV_X1 G3265 (
	 );
   NOR2_X1 G3264 (
	 );
   NAND4_X1 G3263 (
	 );
   NAND3_X1 G3262 (
	 );
   NAND4_X1 G3261 (
	 );
   NAND3_X1 G3260 (
	 );
   NAND4_X1 G3259 (
	 );
   NAND2_X1 G3258 (
	 );
   NOR2_X1 G3257 (
	 );
   INV_X1 G3256 (
	 );
   NOR2_X1 G3255 (
	 );
   NOR2_X1 G3254 (
	 );
   INV_X1 G3253 (
	 );
   NOR2_X1 G3252 (
	 );
   INV_X1 G3251 (
	 );
   MUX2_X1 G3250 (
	 );
   CLKBUF_X1 G3249 (
	 );
   CLKBUF_X1 G3248 (
	 );
   NAND3_X1 G3247 (
	 );
   AOI22_X1 G3246 (
	 );
   AND3_X1 G3245 (
	 );
   NAND2_X1 G3244 (
	 );
   NAND2_X1 G3243 (
	 );
   NAND4_X1 G3242 (
	 );
   NAND3_X1 G3241 (
	 );
   NAND3_X1 G3240 (
	 );
   NAND3_X1 G3239 (
	 );
   NAND2_X1 G3238 (
	 );
   NAND2_X1 G3237 (
	 );
   AND3_X1 G3236 (
	 );
   NAND4_X1 G3235 (
	 );
   NAND4_X1 G3234 (
	 );
   NAND4_X1 G3233 (
	 );
   CLKBUF_X1 G3232 (
	 );
   CLKBUF_X1 G3231 (
	 );
   MUX2_X1 G3230 (
	 );
   CLKBUF_X1 G3229 (
	 );
   MUX2_X1 G3228 (
	 );
   CLKBUF_X1 G3227 (
	 );
   CLKBUF_X1 G3226 (
	 );
   CLKBUF_X1 G3225 (
	 );
   MUX2_X1 G3224 (
	 );
   CLKBUF_X1 G3223 (
	 );
   OAI21_X1 G3222 (
	 );
   NAND3_X1 G3221 (
	 );
   NAND2_X1 G3220 (
	 );
   OAI211_X1 G3219 (
	 );
   XNOR2_X1 G3218 (
	 );
   MUX2_X1 G3217 (
	 );
   CLKBUF_X1 G3216 (
	 );
   NOR2_X1 G3215 (
	 );
   CLKBUF_X1 G3214 (
	 );
   CLKBUF_X1 G3213 (
	 );
   CLKBUF_X1 G3212 (
	 );
   CLKBUF_X1 G3211 (
	 );
   OAI221_X1 G3210 (
	 );
   INV_X1 G3209 (
	 );
   AOI22_X1 G3208 (
	 );
   CLKBUF_X1 G3207 (
	 );
   OAI21_X1 G3206 (
	 );
   INV_X1 G3205 (
	 );
   NOR2_X1 G3204 (
	 );
   NOR2_X1 G3203 (
	 );
   MUX2_X1 G3202 (
	 );
   CLKBUF_X1 G3201 (
	 );
   CLKBUF_X1 G3200 (
	 );
   NOR2_X1 G3199 (
	 );
   INV_X1 G3198 (
	 );
   NAND3_X1 G3197 (
	 );
   CLKBUF_X1 G3196 (
	 );
   CLKBUF_X1 G3195 (
	 );
   MUX2_X1 G3194 (
	 );
   CLKBUF_X1 G3193 (
	 );
   CLKBUF_X1 G3192 (
	 );
   OAI211_X1 G3191 (
	 );
   NAND4_X1 G3190 (
	 );
   NOR3_X1 G3189 (
	 );
   AND3_X1 G3188 (
	 );
   NOR2_X1 G3187 (
	 );
   OAI22_X1 G3186 (
	 );
   INV_X1 G3185 (
	 );
   INV_X1 G3184 (
	 );
   CLKBUF_X1 G3183 (
	 );
   NOR2_X1 G3182 (
	 );
   MUX2_X1 G3181 (
	 );
   OAI21_X1 G3180 (
	 );
   INV_X1 G3179 (
	 );
   AOI22_X1 G3178 (
	 );
   CLKBUF_X1 G3177 (
	 );
   MUX2_X1 G3176 (
	 );
   CLKBUF_X1 G3175 (
	 );
   OAI21_X1 G3174 (
	 );
   INV_X1 G3173 (
	 );
   NAND2_X1 G3172 (
	 );
   OAI22_X1 G3171 (
	 );
   INV_X1 G3170 (
	 );
   CLKBUF_X1 G3169 (
	 );
   CLKBUF_X1 G3168 (
	 );
   MUX2_X1 G3167 (
	 );
   CLKBUF_X1 G3166 (
	 );
   CLKBUF_X1 G3165 (
	 );
   CLKBUF_X1 G3164 (
	 );
   NOR2_X1 G3163 (
	 );
   CLKBUF_X1 G3162 (
	 );
   MUX2_X1 G3161 (
	 );
   CLKBUF_X1 G3160 (
	 );
   CLKBUF_X1 G3159 (
	 );
   CLKBUF_X1 G3158 (
	 );
   CLKBUF_X1 G3157 (
	 );
   AOI21_X1 G3156 (
	 );
   OAI21_X1 G3155 (
	 );
   OAI21_X1 G3154 (
	 );
   NAND2_X1 G3153 (
	 );
   OAI21_X1 G3152 (
	 );
   NAND2_X1 G3151 (
	 );
   CLKBUF_X1 G3150 (
	 );
   CLKBUF_X1 G3149 (
	 );
   CLKBUF_X1 G3148 (
	 );
   NAND3_X1 G3147 (
	 );
   AND3_X1 G3146 (
	 );
   NAND2_X1 G3145 (
	 );
   NAND2_X1 G3144 (
	 );
   NAND2_X1 G3143 (
	 );
   AOI22_X1 G3142 (
	 );
   NAND2_X1 G3141 (
	 );
   AOI22_X1 G3140 (
	 );
   AOI22_X1 G3139 (
	 );
   AND3_X1 G3138 (
	 );
   NAND4_X1 G3137 (
	 );
   NAND4_X1 G3136 (
	 );
   NAND4_X1 G3135 (
	 );
   INV_X1 G3134 (
	 );
   CLKBUF_X1 G3133 (
	 );
   NOR2_X1 G3132 (
	 );
   AND2_X1 G3131 (
	 );
   CLKBUF_X1 G3130 (
	 );
   CLKBUF_X1 G3129 (
	 );
   NAND3_X1 G3128 (
	 );
   NAND4_X1 G3127 (
	 );
   NOR3_X1 G3126 (
	 );
   NAND3_X1 G3125 (
	 );
   NAND4_X1 G3124 (
	 );
   NAND3_X1 G3123 (
	 );
   NAND3_X1 G3122 (
	 );
   OAI22_X1 G3121 (
	 );
   INV_X1 G3120 (
	 );
   AND4_X1 G3119 (
	 );
   NOR2_X1 G3118 (
	 );
   NOR2_X1 G3117 (
	 );
   NOR2_X1 G3116 (
	 );
   NOR4_X1 G3115 (
	 );
   NAND4_X1 G3114 (
	 );
   CLKBUF_X1 G3113 (
	 );
   CLKBUF_X1 G3112 (
	 );
   CLKBUF_X1 G3111 (
	 );
   OAI21_X1 G3110 (
	 );
   INV_X1 G3109 (
	 );
   NAND2_X1 G3108 (
	 );
   CLKBUF_X1 G3107 (
	 );
   OAI21_X1 G3106 (
	 );
   INV_X1 G3105 (
	 );
   NAND2_X1 G3104 (
	 );
   OAI21_X1 G3103 (
	 );
   INV_X1 G3102 (
	 );
   NAND2_X1 G3101 (
	 );
   NAND2_X1 G3100 (
	 );
   AOI22_X1 G3099 (
	 );
   AOI22_X1 G3098 (
	 );
   NAND2_X1 G3097 (
	 );
   AOI22_X1 G3096 (
	 );
   AOI22_X1 G3095 (
	 );
   CLKBUF_X1 G3094 (
	 );
   OAI21_X1 G3093 (
	 );
   INV_X1 G3092 (
	 );
   NAND2_X1 G3091 (
	 );
   CLKBUF_X1 G3090 (
	 );
   CLKBUF_X1 G3089 (
	 );
   CLKBUF_X1 G3088 (
	 );
   MUX2_X1 G3087 (
	 );
   CLKBUF_X1 G3086 (
	 );
   CLKBUF_X1 G3085 (
	 );
   OAI21_X1 G3084 (
	 );
   INV_X1 G3083 (
	 );
   NAND2_X1 G3082 (
	 );
   AOI21_X1 G3081 (
	 );
   OAI21_X1 G3080 (
	 );
   AND2_X1 G3079 (
	 );
   CLKBUF_X1 G3078 (
	 );
   CLKBUF_X1 G3077 (
	 );
   OAI21_X1 G3076 (
	 );
   NAND2_X1 G3075 (
	 );
   OAI221_X1 G3074 (
	 );
   NAND2_X1 G3073 (
	 );
   CLKBUF_X1 G3072 (
	 );
   CLKBUF_X1 G3071 (
	 );
   CLKBUF_X1 G3070 (
	 );
   OAI21_X1 G3069 (
	 );
   INV_X1 G3068 (
	 );
   NAND2_X1 G3067 (
	 );
   CLKBUF_X1 G3066 (
	 );
   OAI21_X1 G3065 (
	 );
   INV_X1 G3064 (
	 );
   NAND2_X1 G3063 (
	 );
   NAND3_X1 G3062 (
	 );
   AOI22_X1 G3061 (
	 );
   AND3_X1 G3060 (
	 );
   NAND2_X1 G3059 (
	 );
   NAND2_X1 G3058 (
	 );
   NAND4_X1 G3057 (
	 );
   NAND3_X1 G3056 (
	 );
   NAND3_X1 G3055 (
	 );
   NAND3_X1 G3054 (
	 );
   NAND2_X1 G3053 (
	 );
   NAND2_X1 G3052 (
	 );
   NAND4_X1 G3051 (
	 );
   NAND3_X1 G3050 (
	 );
   NAND3_X1 G3049 (
	 );
   NAND3_X1 G3048 (
	 );
   NAND2_X1 G3047 (
	 );
   AND3_X1 G3046 (
	 );
   NAND4_X1 G3045 (
	 );
   NAND4_X1 G3044 (
	 );
   NAND4_X1 G3043 (
	 );
   AND2_X1 G3042 (
	 );
   AND2_X1 G3041 (
	 );
   CLKBUF_X1 G3040 (
	 );
   NAND2_X1 G3039 (
	 );
   AOI22_X1 G3038 (
	 );
   AOI22_X1 G3037 (
	 );
   NAND3_X1 G3036 (
	 );
   AOI22_X1 G3035 (
	 );
   AND3_X1 G3034 (
	 );
   NAND2_X1 G3033 (
	 );
   NAND2_X1 G3032 (
	 );
   NAND2_X1 G3031 (
	 );
   AND3_X1 G3030 (
	 );
   NAND4_X1 G3029 (
	 );
   NAND4_X1 G3028 (
	 );
   NAND4_X1 G3027 (
	 );
   OAI21_X1 G3026 (
	 );
   NAND2_X1 G3025 (
	 );
   CLKBUF_X1 G3024 (
	 );
   NOR2_X1 G3023 (
	 );
   INV_X1 G3022 (
	 );
   CLKBUF_X1 G3021 (
	 );
   MUX2_X1 G3020 (
	 );
   CLKBUF_X1 G3019 (
	 );
   NAND4_X1 G3018 (
	 );
   NAND2_X1 G3017 (
	 );
   NAND2_X1 G3016 (
	 );
   AOI22_X1 G3015 (
	 );
   AOI22_X1 G3014 (
	 );
   NAND2_X1 G3013 (
	 );
   NAND2_X1 G3012 (
	 );
   AOI22_X1 G3011 (
	 );
   CLKBUF_X1 G3010 (
	 );
   CLKBUF_X1 G3009 (
	 );
   CLKBUF_X1 G3008 (
	 );
   OAI21_X1 G3007 (
	 );
   INV_X1 G3006 (
	 );
   NAND2_X1 G3005 (
	 );
   NAND2_X1 G3004 (
	 );
   OAI221_X1 G3003 (
	 );
   INV_X1 G3002 (
	 );
   AOI22_X1 G3001 (
	 );
   INV_X1 G3000 (
	 );
   INV_X1 G2999 (
	 );
   AND2_X1 G2998 (
	 );
   CLKBUF_X1 G2997 (
	 );
   AND2_X1 G2996 (
	 );
   OAI21_X1 G2995 (
	 );
   INV_X1 G2994 (
	 );
   NAND2_X1 G2993 (
	 );
   OAI21_X1 G2992 (
	 );
   INV_X1 G2991 (
	 );
   AOI22_X1 G2990 (
	 );
   OAI21_X1 G2989 (
	 );
   INV_X1 G2988 (
	 );
   NAND2_X1 G2987 (
	 );
   NOR2_X1 G2986 (
	 );
   MUX2_X1 G2985 (
	 );
   CLKBUF_X1 G2984 (
	 );
   MUX2_X1 G2983 (
	 );
   CLKBUF_X1 G2982 (
	 );
   CLKBUF_X1 G2981 (
	 );
   CLKBUF_X1 G2980 (
	 );
   OAI21_X1 G2979 (
	 );
   NAND2_X1 G2978 (
	 );
   OAI22_X1 G2977 (
	 );
   CLKBUF_X1 G2976 (
	 );
   CLKBUF_X1 G2975 (
	 );
   AOI21_X1 G2974 (
	 );
   INV_X1 G2973 (
	 );
   NOR2_X1 G2972 (
	 );
   CLKBUF_X1 G2971 (
	 );
   CLKBUF_X1 G2970 (
	 );
   CLKBUF_X1 G2969 (
	 );
   CLKBUF_X1 G2968 (
	 );
   MUX2_X1 G2967 (
	 );
   NOR2_X1 G2966 (
	 );
   OAI21_X1 G2965 (
	 );
   INV_X1 G2964 (
	 );
   NAND2_X1 G2963 (
	 );
   CLKBUF_X1 G2962 (
	 );
   CLKBUF_X1 G2961 (
	 );
   AND2_X1 G2960 (
	 );
   CLKBUF_X1 G2959 (
	 );
   CLKBUF_X1 G2958 (
	 );
   NOR4_X1 G2957 (
	 );
   NAND2_X1 G2956 (
	 );
   INV_X1 G2955 (
	 );
   NAND3_X1 G2954 (
	 );
   INV_X1 G2953 (
	 );
   INV_X1 G2952 (
	 );
   CLKBUF_X1 G2951 (
	 );
   OAI21_X1 G2950 (
	 );
   OAI21_X1 G2949 (
	 );
   NAND2_X1 G2948 (
	 );
   NAND3_X1 G2947 (
	 );
   NOR2_X1 G2946 (
	 );
   NAND3_X1 G2945 (
	 );
   INV_X1 G2944 (
	 );
   NOR2_X1 G2943 (
	 );
   CLKBUF_X1 G2942 (
	 );
   NAND4_X1 G2941 (
	 );
   NAND2_X1 G2940 (
	 );
   NAND2_X1 G2939 (
	 );
   AOI22_X1 G2938 (
	 );
   AOI22_X1 G2937 (
	 );
   NAND2_X1 G2936 (
	 );
   NAND2_X1 G2935 (
	 );
   AOI22_X1 G2934 (
	 );
   OAI21_X1 G2933 (
	 );
   INV_X1 G2932 (
	 );
   NAND2_X1 G2931 (
	 );
   XNOR2_X1 G2930 (
	 );
   NAND2_X1 G2929 (
	 );
   CLKBUF_X1 G2928 (
	 );
   CLKBUF_X1 G2927 (
	 );
   CLKBUF_X1 G2926 (
	 );
   CLKBUF_X1 G2925 (
	 );
   CLKBUF_X1 G2924 (
	 );
   CLKBUF_X1 G2923 (
	 );
   NAND3_X1 G2922 (
	 );
   AOI22_X1 G2921 (
	 );
   AND3_X1 G2920 (
	 );
   NAND2_X1 G2919 (
	 );
   NAND2_X1 G2918 (
	 );
   NAND2_X1 G2917 (
	 );
   AND3_X1 G2916 (
	 );
   NAND4_X1 G2915 (
	 );
   NAND4_X1 G2914 (
	 );
   NAND4_X1 G2913 (
	 );
   CLKBUF_X1 G2912 (
	 );
   MUX2_X1 G2911 (
	 );
   CLKBUF_X1 G2910 (
	 );
   CLKBUF_X1 G2909 (
	 );
   NOR2_X1 G2908 (
	 );
   NAND4_X1 G2907 (
	 );
   NAND2_X1 G2906 (
	 );
   NAND2_X1 G2905 (
	 );
   OAI21_X1 G2904 (
	 );
   NAND3_X1 G2903 (
	 );
   OAI21_X1 G2902 (
	 );
   OAI21_X1 G2901 (
	 );
   XNOR2_X1 G2900 (
	 );
   INV_X1 G2899 (
	 );
   XNOR2_X1 G2898 (
	 );
   NAND3_X1 G2897 (
	 );
   CLKBUF_X1 G2896 (
	 );
   MUX2_X1 G2895 (
	 );
   OAI221_X1 G2894 (
	 );
   AOI22_X1 G2893 (
	 );
   CLKBUF_X1 G2892 (
	 );
   OAI21_X1 G2891 (
	 );
   INV_X1 G2890 (
	 );
   INV_X1 G2889 (
	 );
   INV_X1 G2888 (
	 );
   CLKBUF_X1 G2887 (
	 );
   CLKBUF_X1 G2886 (
	 );
   CLKBUF_X1 G2885 (
	 );
   OAI21_X1 G2884 (
	 );
   INV_X1 G2883 (
	 );
   NAND2_X1 G2882 (
	 );
   OAI221_X1 G2881 (
	 );
   NAND2_X1 G2880 (
	 );
   NAND2_X1 G2879 (
	 );
   AOI22_X1 G2878 (
	 );
   AOI22_X1 G2877 (
	 );
   CLKBUF_X1 G2876 (
	 );
   INV_X1 G2875 (
	 );
   NAND2_X1 G2874 (
	 );
   OAI21_X1 G2873 (
	 );
   INV_X1 G2872 (
	 );
   NAND2_X1 G2871 (
	 );
   CLKBUF_X1 G2870 (
	 );
   CLKBUF_X1 G2869 (
	 );
   CLKBUF_X1 G2868 (
	 );
   CLKBUF_X1 G2867 (
	 );
   CLKBUF_X1 G2866 (
	 );
   OAI21_X1 G2865 (
	 );
   INV_X1 G2864 (
	 );
   NAND2_X1 G2863 (
	 );
   NOR3_X1 G2862 (
	 );
   AOI21_X1 G2861 (
	 );
   AND3_X1 G2860 (
	 );
   CLKBUF_X1 G2859 (
	 );
   AOI21_X1 G2858 (
	 );
   OAI21_X1 G2857 (
	 );
   NAND3_X1 G2856 (
	 );
   OAI21_X1 G2855 (
	 );
   INV_X1 G2854 (
	 );
   INV_X1 G2853 (
	 );
   OAI21_X1 G2852 (
	 );
   INV_X1 G2851 (
	 );
   NAND2_X1 G2850 (
	 );
   CLKBUF_X1 G2849 (
	 );
   MUX2_X1 G2848 (
	 );
   CLKBUF_X1 G2847 (
	 );
   CLKBUF_X1 G2846 (
	 );
   OAI21_X1 G2845 (
	 );
   INV_X1 G2844 (
	 );
   NAND2_X1 G2843 (
	 );
   NAND3_X1 G2842 (
	 );
   NAND2_X1 G2841 (
	 );
   OR2_X1 G2840 (
	 );
   AND4_X1 G2839 (
	 );
   MUX2_X1 G2838 (
	 );
   AND2_X1 G2837 (
	 );
   CLKBUF_X1 G2836 (
	 );
   CLKBUF_X1 G2835 (
	 );
   CLKBUF_X1 G2834 (
	 );
   OAI21_X1 G2833 (
	 );
   INV_X1 G2832 (
	 );
   NAND2_X1 G2831 (
	 );
   OAI21_X1 G2830 (
	 );
   INV_X1 G2829 (
	 );
   AOI22_X1 G2828 (
	 );
   CLKBUF_X1 G2827 (
	 );
   CLKBUF_X1 G2826 (
	 );
   CLKBUF_X1 G2825 (
	 );
   CLKBUF_X1 G2824 (
	 );
   MUX2_X1 G2823 (
	 );
   CLKBUF_X1 G2822 (
	 );
   CLKBUF_X1 G2821 (
	 );
   MUX2_X1 G2820 (
	 );
   CLKBUF_X1 G2819 (
	 );
   CLKBUF_X1 G2818 (
	 );
   AOI21_X1 G2817 (
	 );
   INV_X1 G2816 (
	 );
   CLKBUF_X1 G2815 (
	 );
   CLKBUF_X1 G2814 (
	 );
   CLKBUF_X1 G2813 (
	 );
   NAND2_X1 G2812 (
	 );
   NAND3_X1 G2811 (
	 );
   NAND2_X1 G2810 (
	 );
   INV_X1 G2809 (
	 );
   AOI22_X1 G2808 (
	 );
   AOI22_X1 G2807 (
	 );
   NOR2_X1 G2806 (
	 );
   CLKBUF_X1 G2805 (
	 );
   CLKBUF_X1 G2804 (
	 );
   CLKBUF_X1 G2803 (
	 );
   NAND2_X1 G2802 (
	 );
   AND4_X1 G2801 (
	 );
   NAND2_X1 G2800 (
	 );
   NAND2_X1 G2799 (
	 );
   NAND2_X1 G2798 (
	 );
   NAND2_X1 G2797 (
	 );
   AND4_X1 G2796 (
	 );
   NAND4_X1 G2795 (
	 );
   NAND4_X1 G2794 (
	 );
   NAND3_X1 G2793 (
	 );
   NAND3_X1 G2792 (
	 );
   AND2_X1 G2791 (
	 );
   BUF_X2 G2790 (
	 );
   CLKBUF_X1 G2789 (
	 );
   OAI21_X1 G2788 (
	 );
   INV_X1 G2787 (
	 );
   NAND2_X1 G2786 (
	 );
   CLKBUF_X1 G2785 (
	 );
   CLKBUF_X1 G2784 (
	 );
   CLKBUF_X1 G2783 (
	 );
   CLKBUF_X1 G2782 (
	 );
   CLKBUF_X1 G2781 (
	 );
   MUX2_X1 G2780 (
	 );
   OAI21_X1 G2779 (
	 );
   INV_X1 G2778 (
	 );
   AOI22_X1 G2777 (
	 );
   CLKBUF_X1 G2776 (
	 );
   OAI21_X1 G2775 (
	 );
   INV_X1 G2774 (
	 );
   NAND2_X1 G2773 (
	 );
   OAI21_X1 G2772 (
	 );
   AOI22_X1 G2771 (
	 );
   MUX2_X1 G2770 (
	 );
   NAND2_X1 G2769 (
	 );
   AND4_X1 G2768 (
	 );
   NAND2_X1 G2767 (
	 );
   NAND2_X1 G2766 (
	 );
   NAND2_X1 G2765 (
	 );
   NAND2_X1 G2764 (
	 );
   NAND4_X1 G2763 (
	 );
   NAND3_X1 G2762 (
	 );
   NAND3_X1 G2761 (
	 );
   NAND3_X1 G2760 (
	 );
   NAND2_X1 G2759 (
	 );
   AND4_X1 G2758 (
	 );
   NAND4_X1 G2757 (
	 );
   NAND4_X1 G2756 (
	 );
   NAND3_X1 G2755 (
	 );
   NAND3_X1 G2754 (
	 );
   CLKBUF_X1 G2753 (
	 );
   AOI21_X1 G2752 (
	 );
   INV_X1 G2751 (
	 );
   NOR2_X1 G2750 (
	 );
   NAND2_X1 G2749 (
	 );
   AOI22_X1 G2748 (
	 );
   AOI22_X1 G2747 (
	 );
   CLKBUF_X1 G2746 (
	 );
   CLKBUF_X1 G2745 (
	 );
   CLKBUF_X1 G2744 (
	 );
   MUX2_X1 G2743 (
	 );
   MUX2_X1 G2742 (
	 );
   CLKBUF_X1 G2741 (
	 );
   OAI21_X1 G2740 (
	 );
   INV_X1 G2739 (
	 );
   INV_X1 G2738 (
	 );
   NAND2_X1 G2737 (
	 );
   NOR3_X1 G2736 (
	 );
   INV_X1 G2735 (
	 );
   XNOR2_X1 G2734 (
	 );
   NAND2_X1 G2733 (
	 );
   XNOR2_X1 G2732 (
	 );
   CLKBUF_X1 G2731 (
	 );
   CLKBUF_X1 G2730 (
	 );
   OAI21_X1 G2729 (
	 );
   INV_X1 G2728 (
	 );
   NAND2_X1 G2727 (
	 );
   CLKBUF_X1 G2726 (
	 );
   CLKBUF_X1 G2725 (
	 );
   NAND3_X1 G2724 (
	 );
   AOI22_X1 G2723 (
	 );
   AND3_X1 G2722 (
	 );
   NAND2_X1 G2721 (
	 );
   NAND2_X1 G2720 (
	 );
   NAND2_X1 G2719 (
	 );
   AND3_X1 G2718 (
	 );
   NAND4_X1 G2717 (
	 );
   NAND4_X1 G2716 (
	 );
   NAND4_X1 G2715 (
	 );
   MUX2_X1 G2714 (
	 );
   AOI21_X1 G2713 (
	 );
   NOR2_X1 G2712 (
	 );
   NAND2_X1 G2711 (
	 );
   INV_X1 G2710 (
	 );
   OAI21_X1 G2709 (
	 );
   INV_X1 G2708 (
	 );
   NOR3_X1 G2707 (
	 );
   NAND4_X1 G2706 (
	 );
   INV_X1 G2705 (
	 );
   INV_X1 G2704 (
	 );
   INV_X1 G2703 (
	 );
   CLKBUF_X1 G2702 (
	 );
   CLKBUF_X1 G2701 (
	 );
   CLKBUF_X1 G2700 (
	 );
   OAI221_X1 G2699 (
	 );
   INV_X1 G2698 (
	 );
   INV_X1 G2697 (
	 );
   AOI22_X1 G2696 (
	 );
   CLKBUF_X1 G2695 (
	 );
   CLKBUF_X1 G2694 (
	 );
   CLKBUF_X1 G2693 (
	 );
   AOI21_X1 G2692 (
	 );
   NAND2_X1 G2691 (
	 );
   INV_X1 G2690 (
	 );
   CLKBUF_X1 G2689 (
	 );
   AOI21_X1 G2688 (
	 );
   OAI21_X1 G2687 (
	 );
   NAND2_X1 G2686 (
	 );
   MUX2_X1 G2685 (
	 );
   CLKBUF_X1 G2684 (
	 );
   CLKBUF_X1 G2683 (
	 );
   CLKBUF_X1 G2682 (
	 );
   MUX2_X1 G2681 (
	 );
   CLKBUF_X1 G2680 (
	 );
   CLKBUF_X1 G2679 (
	 );
   CLKBUF_X1 G2678 (
	 );
   CLKBUF_X1 G2677 (
	 );
   MUX2_X1 G2676 (
	 );
   OAI21_X1 G2675 (
	 );
   INV_X1 G2674 (
	 );
   AOI22_X1 G2673 (
	 );
   OAI21_X1 G2672 (
	 );
   INV_X1 G2671 (
	 );
   NAND2_X1 G2670 (
	 );
   CLKBUF_X1 G2669 (
	 );
   CLKBUF_X1 G2668 (
	 );
   CLKBUF_X1 G2667 (
	 );
   CLKBUF_X1 G2666 (
	 );
   CLKBUF_X1 G2665 (
	 );
   AND2_X1 G2664 (
	 );
   INV_X1 G2663 (
	 );
   AOI211_X1 G2662 (
	 );
   INV_X1 G2661 (
	 );
   CLKBUF_X1 G2660 (
	 );
   CLKBUF_X1 G2659 (
	 );
   NOR2_X1 G2658 (
	 );
   AOI21_X1 G2657 (
	 );
   OAI21_X1 G2656 (
	 );
   INV_X1 G2655 (
	 );
   NAND2_X1 G2654 (
	 );
   CLKBUF_X1 G2653 (
	 );
   AOI21_X1 G2652 (
	 );
   INV_X1 G2651 (
	 );
   NAND3_X1 G2650 (
	 );
   AOI21_X1 G2649 (
	 );
   AOI21_X1 G2648 (
	 );
   OAI21_X1 G2647 (
	 );
   INV_X1 G2646 (
	 );
   NOR2_X1 G2645 (
	 );
   INV_X1 G2644 (
	 );
   CLKBUF_X1 G2643 (
	 );
   AOI21_X1 G2642 (
	 );
   INV_X1 G2641 (
	 );
   INV_X1 G2640 (
	 );
   CLKBUF_X1 G2639 (
	 );
   AOI21_X1 G2638 (
	 );
   INV_X1 G2637 (
	 );
   NOR2_X1 G2636 (
	 );
   NOR2_X1 G2635 (
	 );
   CLKBUF_X1 G2634 (
	 );
   CLKBUF_X1 G2633 (
	 );
   CLKBUF_X1 G2632 (
	 );
   OAI211_X1 G2631 (
	 );
   NAND4_X1 G2630 (
	 );
   NOR3_X1 G2629 (
	 );
   AND3_X1 G2628 (
	 );
   NOR2_X1 G2627 (
	 );
   OAI22_X1 G2626 (
	 );
   INV_X1 G2625 (
	 );
   INV_X1 G2624 (
	 );
   NAND2_X1 G2623 (
	 );
   NOR2_X1 G2622 (
	 );
   INV_X1 G2621 (
	 );
   MUX2_X1 G2620 (
	 );
   OAI21_X1 G2619 (
	 );
   INV_X1 G2618 (
	 );
   AOI22_X1 G2617 (
	 );
   OAI21_X1 G2616 (
	 );
   NAND2_X1 G2615 (
	 );
   INV_X1 G2614 (
	 );
   NAND3_X1 G2613 (
	 );
   INV_X1 G2612 (
	 );
   NAND2_X1 G2611 (
	 );
   NAND3_X1 G2610 (
	 );
   INV_X1 G2609 (
	 );
   INV_X1 G2608 (
	 );
   CLKBUF_X1 G2607 (
	 );
   CLKBUF_X1 G2606 (
	 );
   MUX2_X1 G2605 (
	 );
   NAND3_X1 G2604 (
	 );
   AOI22_X1 G2603 (
	 );
   AND3_X1 G2602 (
	 );
   NAND2_X1 G2601 (
	 );
   NAND2_X1 G2600 (
	 );
   NAND2_X1 G2599 (
	 );
   NAND4_X1 G2598 (
	 );
   NAND3_X1 G2597 (
	 );
   NAND3_X1 G2596 (
	 );
   NAND3_X1 G2595 (
	 );
   NAND2_X1 G2594 (
	 );
   AND3_X1 G2593 (
	 );
   NAND4_X1 G2592 (
	 );
   NAND4_X1 G2591 (
	 );
   NAND4_X1 G2590 (
	 );
   NOR2_X1 G2589 (
	 );
   CLKBUF_X1 G2588 (
	 );
   XNOR2_X1 G2587 (
	 );
   NAND2_X1 G2586 (
	 );
   XNOR2_X1 G2585 (
	 );
   CLKBUF_X1 G2584 (
	 );
   CLKBUF_X1 G2583 (
	 );
   NAND2_X1 G2582 (
	 );
   AOI22_X1 G2581 (
	 );
   AOI22_X1 G2580 (
	 );
   OAI21_X1 G2579 (
	 );
   NOR2_X1 G2578 (
	 );
   NOR2_X1 G2577 (
	 );
   INV_X1 G2576 (
	 );
   NOR2_X1 G2575 (
	 );
   INV_X1 G2574 (
	 );
   NAND3_X1 G2573 (
	 );
   MUX2_X1 G2572 (
	 );
   AND2_X1 G2571 (
	 );
   CLKBUF_X1 G2570 (
	 );
   CLKBUF_X1 G2569 (
	 );
   CLKBUF_X1 G2568 (
	 );
   AND2_X1 G2567 (
	 );
   CLKBUF_X1 G2566 (
	 );
   CLKBUF_X1 G2565 (
	 );
   CLKBUF_X1 G2564 (
	 );
   CLKBUF_X1 G2563 (
	 );
   CLKBUF_X1 G2562 (
	 );
   CLKBUF_X1 G2561 (
	 );
   AOI21_X1 G2560 (
	 );
   OAI21_X1 G2559 (
	 );
   NAND2_X1 G2558 (
	 );
   CLKBUF_X1 G2557 (
	 );
   NAND3_X1 G2556 (
	 );
   AND3_X1 G2555 (
	 );
   NAND2_X1 G2554 (
	 );
   NAND2_X1 G2553 (
	 );
   NAND4_X1 G2552 (
	 );
   NAND3_X1 G2551 (
	 );
   NAND3_X1 G2550 (
	 );
   NAND3_X1 G2549 (
	 );
   NAND2_X1 G2548 (
	 );
   NAND2_X1 G2547 (
	 );
   AOI22_X1 G2546 (
	 );
   NAND4_X1 G2545 (
	 );
   NAND3_X1 G2544 (
	 );
   NAND3_X1 G2543 (
	 );
   NAND3_X1 G2542 (
	 );
   NAND2_X1 G2541 (
	 );
   AND3_X1 G2540 (
	 );
   NAND4_X1 G2539 (
	 );
   NAND4_X1 G2538 (
	 );
   NAND4_X1 G2537 (
	 );
   CLKBUF_X1 G2536 (
	 );
   CLKBUF_X1 G2535 (
	 );
   CLKBUF_X1 G2534 (
	 );
   OAI21_X1 G2533 (
	 );
   INV_X1 G2532 (
	 );
   NAND2_X1 G2531 (
	 );
   AND2_X1 G2530 (
	 );
   CLKBUF_X1 G2529 (
	 );
   NAND4_X1 G2528 (
	 );
   AOI22_X1 G2527 (
	 );
   NAND2_X1 G2526 (
	 );
   NOR2_X1 G2525 (
	 );
   NAND2_X1 G2524 (
	 );
   NAND2_X1 G2523 (
	 );
   AOI22_X1 G2522 (
	 );
   AOI22_X1 G2521 (
	 );
   NAND2_X1 G2520 (
	 );
   NAND2_X1 G2519 (
	 );
   AOI22_X1 G2518 (
	 );
   AOI22_X1 G2517 (
	 );
   CLKBUF_X1 G2516 (
	 );
   XNOR2_X1 G2515 (
	 );
   NAND3_X1 G2514 (
	 );
   AND3_X1 G2513 (
	 );
   NAND2_X1 G2512 (
	 );
   NAND2_X1 G2511 (
	 );
   NAND2_X1 G2510 (
	 );
   AOI22_X1 G2509 (
	 );
   NAND4_X1 G2508 (
	 );
   NAND3_X1 G2507 (
	 );
   NAND3_X1 G2506 (
	 );
   NAND3_X1 G2505 (
	 );
   NAND2_X1 G2504 (
	 );
   AND3_X1 G2503 (
	 );
   NAND4_X1 G2502 (
	 );
   NAND4_X1 G2501 (
	 );
   NAND4_X1 G2500 (
	 );
   NAND3_X1 G2499 (
	 );
   OR2_X1 G2498 (
	 );
   NOR3_X1 G2497 (
	 );
   NAND3_X1 G2496 (
	 );
   NAND4_X1 G2495 (
	 );
   NAND3_X1 G2494 (
	 );
   NAND3_X1 G2493 (
	 );
   OAI22_X1 G2492 (
	 );
   INV_X1 G2491 (
	 );
   AND4_X1 G2490 (
	 );
   NOR2_X1 G2489 (
	 );
   NOR2_X1 G2488 (
	 );
   NOR2_X1 G2487 (
	 );
   INV_X1 G2486 (
	 );
   NAND4_X1 G2485 (
	 );
   CLKBUF_X1 G2484 (
	 );
   CLKBUF_X1 G2483 (
	 );
   OAI221_X1 G2482 (
	 );
   INV_X1 G2481 (
	 );
   AOI22_X1 G2480 (
	 );
   CLKBUF_X1 G2479 (
	 );
   NAND2_X1 G2478 (
	 );
   MUX2_X1 G2477 (
	 );
   OAI221_X1 G2476 (
	 );
   INV_X1 G2475 (
	 );
   AOI22_X1 G2474 (
	 );
   BUF_X4 G2473 (
	 );
   CLKBUF_X1 G2472 (
	 );
   CLKBUF_X1 G2471 (
	 );
   CLKBUF_X1 G2470 (
	 );
   CLKBUF_X1 G2469 (
	 );
   MUX2_X1 G2468 (
	 );
   OAI21_X1 G2467 (
	 );
   INV_X1 G2466 (
	 );
   AOI22_X1 G2465 (
	 );
   NAND3_X1 G2464 (
	 );
   AOI22_X1 G2463 (
	 );
   NAND4_X1 G2462 (
	 );
   NAND3_X1 G2461 (
	 );
   NAND3_X1 G2460 (
	 );
   NAND3_X1 G2459 (
	 );
   NAND2_X1 G2458 (
	 );
   AND3_X1 G2457 (
	 );
   NAND2_X1 G2456 (
	 );
   NAND2_X1 G2455 (
	 );
   NAND4_X1 G2454 (
	 );
   NAND3_X1 G2453 (
	 );
   NAND3_X1 G2452 (
	 );
   NAND3_X1 G2451 (
	 );
   NAND2_X1 G2450 (
	 );
   NAND2_X1 G2449 (
	 );
   NAND4_X1 G2448 (
	 );
   NAND3_X1 G2447 (
	 );
   NAND3_X1 G2446 (
	 );
   NAND3_X1 G2445 (
	 );
   NAND2_X1 G2444 (
	 );
   AND3_X1 G2443 (
	 );
   NAND4_X1 G2442 (
	 );
   NAND4_X1 G2441 (
	 );
   NAND4_X1 G2440 (
	 );
   CLKBUF_X1 G2439 (
	 );
   CLKBUF_X1 G2438 (
	 );
   CLKBUF_X1 G2437 (
	 );
   CLKBUF_X1 G2436 (
	 );
   NOR2_X1 G2435 (
	 );
   NOR4_X1 G2434 (
	 );
   NOR2_X1 G2433 (
	 );
   NOR2_X1 G2432 (
	 );
   NAND2_X1 G2431 (
	 );
   NAND2_X1 G2430 (
	 );
   OAI21_X1 G2429 (
	 );
   OAI21_X1 G2428 (
	 );
   XNOR2_X1 G2427 (
	 );
   NAND2_X1 G2426 (
	 );
   XOR2_X1 G2425 (
	 );
   CLKBUF_X1 G2424 (
	 );
   CLKBUF_X1 G2423 (
	 );
   MUX2_X1 G2422 (
	 );
   NOR2_X1 G2421 (
	 );
   NAND3_X1 G2420 (
	 );
   NAND4_X1 G2419 (
	 );
   NOR3_X1 G2418 (
	 );
   NAND3_X1 G2417 (
	 );
   NAND4_X1 G2416 (
	 );
   NAND3_X1 G2415 (
	 );
   NAND3_X1 G2414 (
	 );
   OAI22_X1 G2413 (
	 );
   INV_X1 G2412 (
	 );
   INV_X1 G2411 (
	 );
   AND4_X1 G2410 (
	 );
   NOR2_X1 G2409 (
	 );
   NOR2_X1 G2408 (
	 );
   INV_X1 G2407 (
	 );
   NOR2_X1 G2406 (
	 );
   INV_X1 G2405 (
	 );
   CLKBUF_X1 G2404 (
	 );
   CLKBUF_X1 G2403 (
	 );
   MUX2_X1 G2402 (
	 );
   NOR2_X1 G2401 (
	 );
   CLKBUF_X1 G2400 (
	 );
   AND2_X1 G2399 (
	 );
   NAND4_X1 G2398 (
	 );
   NAND4_X1 G2397 (
	 );
   NAND4_X1 G2396 (
	 );
   NAND4_X1 G2395 (
	 );
   NOR2_X1 G2394 (
	 );
   NAND4_X1 G2393 (
	 );
   NAND4_X1 G2392 (
	 );
   NAND3_X1 G2391 (
	 );
   NAND3_X1 G2390 (
	 );
   NAND4_X1 G2389 (
	 );
   NAND2_X1 G2388 (
	 );
   NAND4_X1 G2387 (
	 );
   NAND4_X1 G2386 (
	 );
   CLKBUF_X1 G2385 (
	 );
   NAND4_X1 G2384 (
	 );
   AOI22_X1 G2383 (
	 );
   NAND2_X1 G2382 (
	 );
   NAND2_X1 G2381 (
	 );
   NAND2_X1 G2380 (
	 );
   NAND4_X1 G2379 (
	 );
   NAND3_X1 G2378 (
	 );
   NAND3_X1 G2377 (
	 );
   NAND3_X1 G2376 (
	 );
   NAND2_X1 G2375 (
	 );
   OAI21_X1 G2374 (
	 );
   INV_X1 G2373 (
	 );
   NAND2_X1 G2372 (
	 );
   CLKBUF_X1 G2371 (
	 );
   CLKBUF_X1 G2370 (
	 );
   NAND3_X1 G2369 (
	 );
   AND3_X1 G2368 (
	 );
   NAND2_X1 G2367 (
	 );
   NAND2_X1 G2366 (
	 );
   NAND4_X1 G2365 (
	 );
   NAND3_X1 G2364 (
	 );
   NAND3_X1 G2363 (
	 );
   NAND3_X1 G2362 (
	 );
   NAND2_X1 G2361 (
	 );
   NAND2_X1 G2360 (
	 );
   NAND4_X1 G2359 (
	 );
   NAND3_X1 G2358 (
	 );
   NAND3_X1 G2357 (
	 );
   NAND3_X1 G2356 (
	 );
   NAND2_X1 G2355 (
	 );
   AOI22_X1 G2354 (
	 );
   AND3_X1 G2353 (
	 );
   NAND4_X1 G2352 (
	 );
   NAND4_X1 G2351 (
	 );
   NAND4_X1 G2350 (
	 );
   CLKBUF_X1 G2349 (
	 );
   AND2_X1 G2348 (
	 );
   CLKBUF_X1 G2347 (
	 );
   NOR2_X1 G2346 (
	 );
   CLKBUF_X1 G2345 (
	 );
   NAND3_X1 G2344 (
	 );
   AOI22_X1 G2343 (
	 );
   AND3_X1 G2342 (
	 );
   NAND2_X1 G2341 (
	 );
   NAND2_X1 G2340 (
	 );
   NAND2_X1 G2339 (
	 );
   AND3_X1 G2338 (
	 );
   NAND4_X1 G2337 (
	 );
   NAND4_X1 G2336 (
	 );
   NAND4_X1 G2335 (
	 );
   MUX2_X1 G2334 (
	 );
   CLKBUF_X1 G2333 (
	 );
   MUX2_X1 G2332 (
	 );
   CLKBUF_X1 G2331 (
	 );
   CLKBUF_X1 G2330 (
	 );
   NAND3_X1 G2329 (
	 );
   AOI22_X1 G2328 (
	 );
   NAND4_X1 G2327 (
	 );
   NAND3_X1 G2326 (
	 );
   NAND3_X1 G2325 (
	 );
   NAND3_X1 G2324 (
	 );
   NAND2_X1 G2323 (
	 );
   AND3_X1 G2322 (
	 );
   NAND2_X1 G2321 (
	 );
   NAND2_X1 G2320 (
	 );
   NAND2_X1 G2319 (
	 );
   AND3_X1 G2318 (
	 );
   NAND4_X1 G2317 (
	 );
   NAND4_X1 G2316 (
	 );
   NAND4_X1 G2315 (
	 );
   CLKBUF_X1 G2314 (
	 );
   NOR3_X1 G2313 (
	 );
   INV_X1 G2312 (
	 );
   CLKBUF_X1 G2311 (
	 );
   OAI21_X1 G2310 (
	 );
   INV_X1 G2309 (
	 );
   NAND2_X1 G2308 (
	 );
   OAI21_X1 G2307 (
	 );
   INV_X1 G2306 (
	 );
   AOI22_X1 G2305 (
	 );
   NAND4_X1 G2304 (
	 );
   AOI22_X1 G2303 (
	 );
   NAND4_X1 G2302 (
	 );
   NAND3_X1 G2301 (
	 );
   NAND3_X1 G2300 (
	 );
   NAND3_X1 G2299 (
	 );
   NAND2_X1 G2298 (
	 );
   NAND2_X1 G2297 (
	 );
   NAND2_X1 G2296 (
	 );
   NAND4_X1 G2295 (
	 );
   NAND3_X1 G2294 (
	 );
   NAND3_X1 G2293 (
	 );
   NAND3_X1 G2292 (
	 );
   NAND2_X1 G2291 (
	 );
   NAND2_X1 G2290 (
	 );
   OAI21_X1 G2289 (
	 );
   INV_X1 G2288 (
	 );
   NAND2_X1 G2287 (
	 );
   CLKBUF_X1 G2286 (
	 );
   OAI221_X1 G2285 (
	 );
   INV_X1 G2284 (
	 );
   INV_X1 G2283 (
	 );
   AOI22_X1 G2282 (
	 );
   CLKBUF_X1 G2281 (
	 );
   AOI21_X1 G2280 (
	 );
   INV_X1 G2279 (
	 );
   NOR2_X1 G2278 (
	 );
   NOR2_X1 G2277 (
	 );
   CLKBUF_X1 G2276 (
	 );
   CLKBUF_X1 G2275 (
	 );
   OAI21_X1 G2274 (
	 );
   NAND2_X1 G2273 (
	 );
   OAI221_X1 G2272 (
	 );
   NAND2_X1 G2271 (
	 );
   CLKBUF_X1 G2270 (
	 );
   CLKBUF_X1 G2269 (
	 );
   OAI21_X1 G2268 (
	 );
   INV_X1 G2267 (
	 );
   NAND2_X1 G2266 (
	 );
   NAND2_X1 G2265 (
	 );
   CLKBUF_X1 G2264 (
	 );
   CLKBUF_X1 G2263 (
	 );
   OAI21_X1 G2262 (
	 );
   INV_X1 G2261 (
	 );
   NAND2_X1 G2260 (
	 );
   CLKBUF_X1 G2259 (
	 );
   MUX2_X1 G2258 (
	 );
   CLKBUF_X1 G2257 (
	 );
   OAI21_X1 G2256 (
	 );
   INV_X1 G2255 (
	 );
   NAND2_X1 G2254 (
	 );
   CLKBUF_X1 G2253 (
	 );
   AND2_X1 G2252 (
	 );
   CLKBUF_X1 G2251 (
	 );
   CLKBUF_X1 G2250 (
	 );
   CLKBUF_X1 G2249 (
	 );
   CLKBUF_X1 G2248 (
	 );
   CLKBUF_X1 G2247 (
	 );
   MUX2_X1 G2246 (
	 );
   AND2_X1 G2245 (
	 );
   NOR2_X1 G2244 (
	 );
   NOR3_X1 G2243 (
	 );
   NOR3_X1 G2242 (
	 );
   CLKBUF_X1 G2241 (
	 );
   NAND2_X1 G2240 (
	 );
   AOI22_X1 G2239 (
	 );
   AOI22_X1 G2238 (
	 );
   CLKBUF_X1 G2237 (
	 );
   CLKBUF_X1 G2236 (
	 );
   OAI221_X1 G2235 (
	 );
   INV_X1 G2234 (
	 );
   INV_X1 G2233 (
	 );
   AOI22_X1 G2232 (
	 );
   CLKBUF_X1 G2231 (
	 );
   NOR2_X1 G2230 (
	 );
   XNOR2_X1 G2229 (
	 );
   NAND2_X1 G2228 (
	 );
   XNOR2_X1 G2227 (
	 );
   XNOR2_X1 G2226 (
	 );
   CLKBUF_X1 G2225 (
	 );
   MUX2_X1 G2224 (
	 );
   MUX2_X1 G2223 (
	 );
   CLKBUF_X1 G2222 (
	 );
   CLKBUF_X1 G2221 (
	 );
   CLKBUF_X1 G2220 (
	 );
   OAI221_X1 G2219 (
	 );
   INV_X1 G2218 (
	 );
   AOI22_X1 G2217 (
	 );
   OAI21_X1 G2216 (
	 );
   INV_X1 G2215 (
	 );
   NAND2_X1 G2214 (
	 );
   AND2_X1 G2213 (
	 );
   INV_X1 G2212 (
	 );
   NAND4_X1 G2211 (
	 );
   AOI22_X1 G2210 (
	 );
   NAND4_X1 G2209 (
	 );
   NAND3_X1 G2208 (
	 );
   NAND3_X1 G2207 (
	 );
   NAND3_X1 G2206 (
	 );
   NAND2_X1 G2205 (
	 );
   NAND2_X1 G2204 (
	 );
   NAND4_X1 G2203 (
	 );
   NAND3_X1 G2202 (
	 );
   NAND3_X1 G2201 (
	 );
   NAND3_X1 G2200 (
	 );
   NAND2_X1 G2199 (
	 );
   NAND2_X1 G2198 (
	 );
   NAND2_X1 G2197 (
	 );
   OAI21_X1 G2196 (
	 );
   OAI21_X1 G2195 (
	 );
   NOR2_X1 G2194 (
	 );
   INV_X1 G2193 (
	 );
   NOR2_X1 G2192 (
	 );
   INV_X1 G2191 (
	 );
   NAND2_X1 G2190 (
	 );
   INV_X1 G2189 (
	 );
   CLKBUF_X1 G2188 (
	 );
   NOR3_X1 G2187 (
	 );
   AOI21_X1 G2186 (
	 );
   AND3_X1 G2185 (
	 );
   AOI21_X1 G2184 (
	 );
   INV_X1 G2183 (
	 );
   NOR3_X1 G2182 (
	 );
   INV_X1 G2181 (
	 );
   NOR2_X1 G2180 (
	 );
   NOR3_X1 G2179 (
	 );
   NOR2_X1 G2178 (
	 );
   NOR3_X1 G2177 (
	 );
   XNOR2_X1 G2176 (
	 );
   NAND2_X1 G2175 (
	 );
   CLKBUF_X1 G2174 (
	 );
   CLKBUF_X1 G2173 (
	 );
   CLKBUF_X1 G2172 (
	 );
   NOR2_X1 G2171 (
	 );
   MUX2_X1 G2170 (
	 );
   OAI21_X1 G2169 (
	 );
   INV_X1 G2168 (
	 );
   AOI22_X1 G2167 (
	 );
   NOR2_X1 G2166 (
	 );
   CLKBUF_X1 G2165 (
	 );
   CLKBUF_X1 G2164 (
	 );
   CLKBUF_X1 G2163 (
	 );
   AND2_X1 G2162 (
	 );
   CLKBUF_X1 G2161 (
	 );
   CLKBUF_X1 G2160 (
	 );
   NAND4_X1 G2159 (
	 );
   NAND4_X1 G2158 (
	 );
   OR2_X1 G2157 (
	 );
   OR2_X1 G2156 (
	 );
   INV_X1 G2155 (
	 );
   NOR2_X1 G2154 (
	 );
   AND2_X1 G2153 (
	 );
   NAND4_X1 G2152 (
	 );
   NAND4_X1 G2151 (
	 );
   NAND3_X1 G2150 (
	 );
   NAND3_X1 G2149 (
	 );
   NAND4_X1 G2148 (
	 );
   NOR2_X1 G2147 (
	 );
   CLKBUF_X1 G2146 (
	 );
   NOR2_X1 G2145 (
	 );
   AOI21_X1 G2144 (
	 );
   INV_X1 G2143 (
	 );
   INV_X1 G2142 (
	 );
   CLKBUF_X1 G2141 (
	 );
   MUX2_X1 G2140 (
	 );
   CLKBUF_X1 G2139 (
	 );
   CLKBUF_X1 G2138 (
	 );
   CLKBUF_X1 G2137 (
	 );
   CLKBUF_X1 G2136 (
	 );
   CLKBUF_X1 G2135 (
	 );
   CLKBUF_X1 G2134 (
	 );
   CLKBUF_X1 G2133 (
	 );
   OAI21_X1 G2132 (
	 );
   INV_X1 G2131 (
	 );
   NAND2_X1 G2130 (
	 );
   OAI21_X1 G2129 (
	 );
   INV_X1 G2128 (
	 );
   AOI22_X1 G2127 (
	 );
   AND2_X1 G2126 (
	 );
   OAI21_X1 G2125 (
	 );
   INV_X1 G2124 (
	 );
   NAND2_X1 G2123 (
	 );
   OAI221_X1 G2122 (
	 );
   NAND2_X1 G2121 (
	 );
   CLKBUF_X1 G2120 (
	 );
   OAI21_X1 G2119 (
	 );
   NAND2_X1 G2118 (
	 );
   NAND3_X1 G2117 (
	 );
   AOI22_X1 G2116 (
	 );
   NAND4_X1 G2115 (
	 );
   NAND3_X1 G2114 (
	 );
   NAND3_X1 G2113 (
	 );
   NAND3_X1 G2112 (
	 );
   NAND2_X1 G2111 (
	 );
   AND3_X1 G2110 (
	 );
   NAND2_X1 G2109 (
	 );
   NAND2_X1 G2108 (
	 );
   NAND4_X1 G2107 (
	 );
   NAND3_X1 G2106 (
	 );
   NAND3_X1 G2105 (
	 );
   NAND3_X1 G2104 (
	 );
   NAND2_X1 G2103 (
	 );
   NAND2_X1 G2102 (
	 );
   AND3_X1 G2101 (
	 );
   NAND4_X1 G2100 (
	 );
   NAND4_X1 G2099 (
	 );
   NAND4_X1 G2098 (
	 );
   CLKBUF_X1 G2097 (
	 );
   CLKBUF_X1 G2096 (
	 );
   CLKBUF_X1 G2095 (
	 );
   CLKBUF_X1 G2094 (
	 );
   NAND2_X1 G2093 (
	 );
   AOI22_X1 G2092 (
	 );
   AOI22_X1 G2091 (
	 );
   CLKBUF_X1 G2090 (
	 );
   CLKBUF_X1 G2089 (
	 );
   NAND2_X1 G2088 (
	 );
   AOI22_X1 G2087 (
	 );
   AOI22_X1 G2086 (
	 );
   CLKBUF_X1 G2085 (
	 );
   CLKBUF_X1 G2084 (
	 );
   AND2_X1 G2083 (
	 );
   CLKBUF_X1 G2082 (
	 );
   XNOR2_X1 G2081 (
	 );
   XNOR2_X1 G2080 (
	 );
   MUX2_X1 G2079 (
	 );
   CLKBUF_X1 G2078 (
	 );
   CLKBUF_X1 G2077 (
	 );
   NAND3_X1 G2076 (
	 );
   AOI22_X1 G2075 (
	 );
   AND3_X1 G2074 (
	 );
   NAND2_X1 G2073 (
	 );
   NAND2_X1 G2072 (
	 );
   NAND2_X1 G2071 (
	 );
   NAND4_X1 G2070 (
	 );
   NAND3_X1 G2069 (
	 );
   NAND3_X1 G2068 (
	 );
   NAND3_X1 G2067 (
	 );
   NAND2_X1 G2066 (
	 );
   AND3_X1 G2065 (
	 );
   NAND4_X1 G2064 (
	 );
   NAND4_X1 G2063 (
	 );
   NAND4_X1 G2062 (
	 );
   OAI221_X1 G2061 (
	 );
   INV_X1 G2060 (
	 );
   INV_X1 G2059 (
	 );
   AOI22_X1 G2058 (
	 );
   CLKBUF_X1 G2057 (
	 );
   CLKBUF_X1 G2056 (
	 );
   CLKBUF_X1 G2055 (
	 );
   CLKBUF_X1 G2054 (
	 );
   OAI21_X1 G2053 (
	 );
   INV_X1 G2052 (
	 );
   NAND2_X1 G2051 (
	 );
   OAI21_X1 G2050 (
	 );
   INV_X1 G2049 (
	 );
   AOI22_X1 G2048 (
	 );
   CLKBUF_X1 G2047 (
	 );
   MUX2_X1 G2046 (
	 );
   NAND2_X1 G2045 (
	 );
   AOI22_X1 G2044 (
	 );
   AOI22_X1 G2043 (
	 );
   MUX2_X1 G2042 (
	 );
   CLKBUF_X1 G2041 (
	 );
   CLKBUF_X1 G2040 (
	 );
   CLKBUF_X1 G2039 (
	 );
   NAND2_X1 G2038 (
	 );
   INV_X1 G2037 (
	 );
   OAI21_X1 G2036 (
	 );
   NOR2_X1 G2035 (
	 );
   INV_X1 G2034 (
	 );
   CLKBUF_X1 G2033 (
	 );
   AND2_X1 G2032 (
	 );
   INV_X1 G2031 (
	 );
   AOI211_X1 G2030 (
	 );
   AOI21_X1 G2029 (
	 );
   OAI21_X1 G2028 (
	 );
   INV_X1 G2027 (
	 );
   NOR2_X1 G2026 (
	 );
   INV_X1 G2025 (
	 );
   INV_X1 G2024 (
	 );
   INV_X1 G2023 (
	 );
   CLKBUF_X1 G2022 (
	 );
   CLKBUF_X1 G2021 (
	 );
   CLKBUF_X1 G2020 (
	 );
   CLKBUF_X1 G2019 (
	 );
   NAND2_X1 G2018 (
	 );
   AND4_X1 G2017 (
	 );
   NAND2_X1 G2016 (
	 );
   NAND2_X1 G2015 (
	 );
   NAND4_X1 G2014 (
	 );
   NAND3_X1 G2013 (
	 );
   NAND3_X1 G2012 (
	 );
   NAND3_X1 G2011 (
	 );
   NAND2_X1 G2010 (
	 );
   NAND2_X1 G2009 (
	 );
   NAND4_X1 G2008 (
	 );
   NAND3_X1 G2007 (
	 );
   NAND3_X1 G2006 (
	 );
   NAND3_X1 G2005 (
	 );
   NAND2_X1 G2004 (
	 );
   NAND2_X1 G2003 (
	 );
   NAND4_X1 G2002 (
	 );
   NAND3_X1 G2001 (
	 );
   NAND3_X1 G2000 (
	 );
   NAND3_X1 G1999 (
	 );
   NAND2_X1 G1998 (
	 );
   AND4_X1 G1997 (
	 );
   NAND4_X1 G1996 (
	 );
   NAND4_X1 G1995 (
	 );
   NAND3_X1 G1994 (
	 );
   NAND3_X1 G1993 (
	 );
   CLKBUF_X1 G1992 (
	 );
   CLKBUF_X1 G1991 (
	 );
   OAI221_X1 G1990 (
	 );
   INV_X1 G1989 (
	 );
   INV_X1 G1988 (
	 );
   AOI22_X1 G1987 (
	 );
   CLKBUF_X1 G1986 (
	 );
   CLKBUF_X1 G1985 (
	 );
   NAND2_X1 G1984 (
	 );
   AOI22_X1 G1983 (
	 );
   AOI22_X1 G1982 (
	 );
   AND2_X1 G1981 (
	 );
   CLKBUF_X1 G1980 (
	 );
   CLKBUF_X1 G1979 (
	 );
   CLKBUF_X1 G1978 (
	 );
   CLKBUF_X1 G1977 (
	 );
   CLKBUF_X1 G1976 (
	 );
   CLKBUF_X1 G1975 (
	 );
   CLKBUF_X1 G1974 (
	 );
   CLKBUF_X1 G1973 (
	 );
   CLKBUF_X1 G1972 (
	 );
   NOR2_X1 G1971 (
	 );
   INV_X1 G1970 (
	 );
   NOR2_X1 G1969 (
	 );
   NAND2_X1 G1968 (
	 );
   OAI221_X1 G1967 (
	 );
   INV_X1 G1966 (
	 );
   AOI22_X1 G1965 (
	 );
   BUF_X4 G1964 (
	 );
   OAI221_X1 G1963 (
	 );
   INV_X1 G1962 (
	 );
   INV_X1 G1961 (
	 );
   AOI22_X1 G1960 (
	 );
   CLKBUF_X1 G1959 (
	 );
   MUX2_X1 G1958 (
	 );
   OAI21_X1 G1957 (
	 );
   INV_X1 G1956 (
	 );
   AOI22_X1 G1955 (
	 );
   CLKBUF_X1 G1954 (
	 );
   CLKBUF_X1 G1953 (
	 );
   OAI21_X1 G1952 (
	 );
   INV_X1 G1951 (
	 );
   NAND2_X1 G1950 (
	 );
   OAI221_X1 G1949 (
	 );
   INV_X1 G1948 (
	 );
   NAND2_X1 G1947 (
	 );
   NOR2_X1 G1946 (
	 );
   BUF_X4 G1945 (
	 );
   CLKBUF_X1 G1944 (
	 );
   CLKBUF_X1 G1943 (
	 );
   NAND3_X1 G1942 (
	 );
   AOI22_X1 G1941 (
	 );
   NAND4_X1 G1940 (
	 );
   NAND3_X1 G1939 (
	 );
   NAND3_X1 G1938 (
	 );
   NAND3_X1 G1937 (
	 );
   NAND2_X1 G1936 (
	 );
   AND3_X1 G1935 (
	 );
   NAND2_X1 G1934 (
	 );
   NAND2_X1 G1933 (
	 );
   NAND4_X1 G1932 (
	 );
   NAND3_X1 G1931 (
	 );
   NAND3_X1 G1930 (
	 );
   NAND3_X1 G1929 (
	 );
   NAND2_X1 G1928 (
	 );
   NAND2_X1 G1927 (
	 );
   NAND4_X1 G1926 (
	 );
   NAND3_X1 G1925 (
	 );
   NAND3_X1 G1924 (
	 );
   NAND3_X1 G1923 (
	 );
   NAND2_X1 G1922 (
	 );
   AND3_X1 G1921 (
	 );
   NAND4_X1 G1920 (
	 );
   NAND4_X1 G1919 (
	 );
   NAND4_X1 G1918 (
	 );
   OAI21_X1 G1917 (
	 );
   INV_X1 G1916 (
	 );
   NAND2_X1 G1915 (
	 );
   OAI221_X1 G1914 (
	 );
   INV_X1 G1913 (
	 );
   INV_X1 G1912 (
	 );
   AOI22_X1 G1911 (
	 );
   CLKBUF_X1 G1910 (
	 );
   AOI21_X1 G1909 (
	 );
   NAND2_X1 G1908 (
	 );
   AOI22_X1 G1907 (
	 );
   AOI22_X1 G1906 (
	 );
   MUX2_X1 G1905 (
	 );
   AND2_X1 G1904 (
	 );
   CLKBUF_X1 G1903 (
	 );
   CLKBUF_X1 G1902 (
	 );
   CLKBUF_X1 G1901 (
	 );
   NAND2_X1 G1900 (
	 );
   AOI22_X1 G1899 (
	 );
   AOI22_X1 G1898 (
	 );
   OAI21_X1 G1897 (
	 );
   INV_X1 G1896 (
	 );
   NAND2_X1 G1895 (
	 );
   CLKBUF_X1 G1894 (
	 );
   NAND2_X1 G1893 (
	 );
   AND4_X1 G1892 (
	 );
   NAND2_X1 G1891 (
	 );
   NAND2_X1 G1890 (
	 );
   NAND2_X1 G1889 (
	 );
   NAND2_X1 G1888 (
	 );
   NAND4_X1 G1887 (
	 );
   NAND3_X1 G1886 (
	 );
   NAND3_X1 G1885 (
	 );
   NAND3_X1 G1884 (
	 );
   NAND2_X1 G1883 (
	 );
   AND4_X1 G1882 (
	 );
   NAND4_X1 G1881 (
	 );
   NAND4_X1 G1880 (
	 );
   NAND3_X1 G1879 (
	 );
   NAND3_X1 G1878 (
	 );
   CLKBUF_X1 G1877 (
	 );
   CLKBUF_X1 G1876 (
	 );
   MUX2_X1 G1875 (
	 );
   CLKBUF_X1 G1874 (
	 );
   CLKBUF_X1 G1873 (
	 );
   NOR2_X1 G1872 (
	 );
   XNOR2_X1 G1871 (
	 );
   INV_X1 G1870 (
	 );
   NAND4_X1 G1869 (
	 );
   NAND2_X1 G1868 (
	 );
   OR2_X1 G1867 (
	 );
   OAI21_X1 G1866 (
	 );
   XNOR2_X1 G1865 (
	 );
   OR2_X1 G1864 (
	 );
   NAND2_X1 G1863 (
	 );
   OAI21_X1 G1862 (
	 );
   INV_X1 G1861 (
	 );
   CLKBUF_X1 G1860 (
	 );
   MUX2_X1 G1859 (
	 );
   AOI21_X1 G1858 (
	 );
   INV_X1 G1857 (
	 );
   NOR2_X1 G1856 (
	 );
   CLKBUF_X1 G1855 (
	 );
   CLKBUF_X1 G1854 (
	 );
   CLKBUF_X1 G1853 (
	 );
   NAND3_X1 G1852 (
	 );
   NAND4_X1 G1851 (
	 );
   NOR3_X1 G1850 (
	 );
   NAND3_X1 G1849 (
	 );
   NAND4_X1 G1848 (
	 );
   NAND3_X1 G1847 (
	 );
   NAND3_X1 G1846 (
	 );
   OAI22_X1 G1845 (
	 );
   INV_X1 G1844 (
	 );
   AND4_X1 G1843 (
	 );
   NOR2_X1 G1842 (
	 );
   NOR2_X1 G1841 (
	 );
   INV_X1 G1840 (
	 );
   NOR2_X1 G1839 (
	 );
   INV_X1 G1838 (
	 );
   OAI21_X1 G1837 (
	 );
   INV_X1 G1836 (
	 );
   NAND2_X1 G1835 (
	 );
   AND2_X1 G1834 (
	 );
   CLKBUF_X1 G1833 (
	 );
   OAI221_X1 G1832 (
	 );
   INV_X1 G1831 (
	 );
   INV_X1 G1830 (
	 );
   AOI22_X1 G1829 (
	 );
   CLKBUF_X1 G1828 (
	 );
   NAND4_X1 G1827 (
	 );
   NAND2_X1 G1826 (
	 );
   NAND2_X1 G1825 (
	 );
   NAND2_X1 G1824 (
	 );
   NAND4_X1 G1823 (
	 );
   NAND3_X1 G1822 (
	 );
   NAND3_X1 G1821 (
	 );
   NAND3_X1 G1820 (
	 );
   NAND2_X1 G1819 (
	 );
   AOI22_X1 G1818 (
	 );
   NAND2_X1 G1817 (
	 );
   AOI22_X1 G1816 (
	 );
   AOI22_X1 G1815 (
	 );
   NOR2_X1 G1814 (
	 );
   BUF_X4 G1813 (
	 );
   AOI21_X1 G1812 (
	 );
   INV_X1 G1811 (
	 );
   INV_X1 G1810 (
	 );
   CLKBUF_X1 G1809 (
	 );
   CLKBUF_X1 G1808 (
	 );
   NAND3_X1 G1807 (
	 );
   AOI22_X1 G1806 (
	 );
   NAND4_X1 G1805 (
	 );
   NAND3_X1 G1804 (
	 );
   NAND3_X1 G1803 (
	 );
   NAND3_X1 G1802 (
	 );
   NAND2_X1 G1801 (
	 );
   AND3_X1 G1800 (
	 );
   NAND2_X1 G1799 (
	 );
   NAND2_X1 G1798 (
	 );
   NAND4_X1 G1797 (
	 );
   NAND3_X1 G1796 (
	 );
   NAND3_X1 G1795 (
	 );
   NAND3_X1 G1794 (
	 );
   NAND2_X1 G1793 (
	 );
   NAND2_X1 G1792 (
	 );
   NAND4_X1 G1791 (
	 );
   NAND3_X1 G1790 (
	 );
   NAND3_X1 G1789 (
	 );
   NAND3_X1 G1788 (
	 );
   NAND2_X1 G1787 (
	 );
   AND3_X1 G1786 (
	 );
   NAND4_X1 G1785 (
	 );
   NAND4_X1 G1784 (
	 );
   NAND4_X1 G1783 (
	 );
   CLKBUF_X1 G1782 (
	 );
   CLKBUF_X1 G1781 (
	 );
   CLKBUF_X1 G1780 (
	 );
   CLKBUF_X1 G1779 (
	 );
   CLKBUF_X1 G1778 (
	 );
   CLKBUF_X1 G1777 (
	 );
   AOI21_X1 G1776 (
	 );
   INV_X1 G1775 (
	 );
   NAND3_X1 G1774 (
	 );
   AOI22_X1 G1773 (
	 );
   NAND4_X1 G1772 (
	 );
   NAND3_X1 G1771 (
	 );
   NAND3_X1 G1770 (
	 );
   NAND3_X1 G1769 (
	 );
   NAND2_X1 G1768 (
	 );
   AND3_X1 G1767 (
	 );
   NAND2_X1 G1766 (
	 );
   NAND2_X1 G1765 (
	 );
   NAND4_X1 G1764 (
	 );
   NAND3_X1 G1763 (
	 );
   NAND3_X1 G1762 (
	 );
   NAND3_X1 G1761 (
	 );
   NAND2_X1 G1760 (
	 );
   NAND2_X1 G1759 (
	 );
   NAND4_X1 G1758 (
	 );
   NAND3_X1 G1757 (
	 );
   NAND3_X1 G1756 (
	 );
   NAND3_X1 G1755 (
	 );
   NAND2_X1 G1754 (
	 );
   AND3_X1 G1753 (
	 );
   NAND4_X1 G1752 (
	 );
   NAND4_X1 G1751 (
	 );
   NAND4_X1 G1750 (
	 );
   CLKBUF_X1 G1749 (
	 );
   CLKBUF_X1 G1748 (
	 );
   CLKBUF_X1 G1747 (
	 );
   MUX2_X1 G1746 (
	 );
   OAI21_X1 G1745 (
	 );
   INV_X1 G1744 (
	 );
   AOI22_X1 G1743 (
	 );
   CLKBUF_X1 G1742 (
	 );
   AND2_X1 G1741 (
	 );
   NAND2_X1 G1740 (
	 );
   INV_X1 G1739 (
	 );
   NAND2_X1 G1738 (
	 );
   CLKBUF_X1 G1737 (
	 );
   CLKBUF_X1 G1736 (
	 );
   CLKBUF_X1 G1735 (
	 );
   AOI21_X1 G1734 (
	 );
   INV_X1 G1733 (
	 );
   NAND3_X1 G1732 (
	 );
   AOI22_X1 G1731 (
	 );
   AND3_X1 G1730 (
	 );
   NAND2_X1 G1729 (
	 );
   NAND2_X1 G1728 (
	 );
   NAND4_X1 G1727 (
	 );
   NAND3_X1 G1726 (
	 );
   NAND3_X1 G1725 (
	 );
   NAND3_X1 G1724 (
	 );
   NAND2_X1 G1723 (
	 );
   NAND2_X1 G1722 (
	 );
   NAND4_X1 G1721 (
	 );
   NAND3_X1 G1720 (
	 );
   NAND3_X1 G1719 (
	 );
   NAND3_X1 G1718 (
	 );
   NAND2_X1 G1717 (
	 );
   AND3_X1 G1716 (
	 );
   NAND4_X1 G1715 (
	 );
   NAND4_X1 G1714 (
	 );
   NAND4_X1 G1713 (
	 );
   INV_X1 G1712 (
	 );
   NAND2_X1 G1711 (
	 );
   NAND2_X1 G1710 (
	 );
   INV_X1 G1709 (
	 );
   NAND2_X1 G1708 (
	 );
   OAI21_X1 G1707 (
	 );
   INV_X1 G1706 (
	 );
   NAND2_X1 G1705 (
	 );
   AND2_X1 G1704 (
	 );
   XOR2_X1 G1703 (
	 );
   NAND3_X1 G1702 (
	 );
   NAND4_X1 G1701 (
	 );
   NOR3_X1 G1700 (
	 );
   NAND3_X1 G1699 (
	 );
   NAND4_X1 G1698 (
	 );
   NAND3_X1 G1697 (
	 );
   NAND3_X1 G1696 (
	 );
   OAI22_X1 G1695 (
	 );
   INV_X1 G1694 (
	 );
   INV_X1 G1693 (
	 );
   AND4_X1 G1692 (
	 );
   NOR2_X1 G1691 (
	 );
   NOR2_X1 G1690 (
	 );
   INV_X1 G1689 (
	 );
   NOR2_X1 G1688 (
	 );
   AOI21_X1 G1687 (
	 );
   INV_X1 G1686 (
	 );
   INV_X1 G1685 (
	 );
   NOR3_X1 G1684 (
	 );
   NOR2_X1 G1683 (
	 );
   XNOR2_X1 G1682 (
	 );
   NAND2_X1 G1681 (
	 );
   XNOR2_X1 G1680 (
	 );
   XNOR2_X1 G1679 (
	 );
   NAND2_X1 G1678 (
	 );
   NAND3_X1 G1677 (
	 );
   NAND2_X1 G1676 (
	 );
   INV_X1 G1675 (
	 );
   NOR2_X1 G1674 (
	 );
   AOI22_X1 G1673 (
	 );
   AOI22_X1 G1672 (
	 );
   NOR2_X1 G1671 (
	 );
   INV_X1 G1670 (
	 );
   AND2_X1 G1669 (
	 );
   CLKBUF_X1 G1668 (
	 );
   OAI21_X1 G1667 (
	 );
   NAND2_X1 G1666 (
	 );
   INV_X1 G1665 (
	 );
   NOR2_X1 G1664 (
	 );
   XNOR2_X1 G1663 (
	 );
   OR4_X1 G1662 (
	 );
   NOR2_X1 G1661 (
	 );
   AND2_X1 G1660 (
	 );
   NOR2_X1 G1659 (
	 );
   NOR2_X1 G1658 (
	 );
   INV_X1 G1657 (
	 );
   NAND3_X1 G1656 (
	 );
   CLKBUF_X1 G1655 (
	 );
   OAI221_X1 G1654 (
	 );
   NAND2_X1 G1653 (
	 );
   NAND2_X1 G1652 (
	 );
   NAND2_X1 G1651 (
	 );
   OAI21_X1 G1650 (
	 );
   NOR2_X1 G1649 (
	 );
   NAND3_X1 G1648 (
	 );
   AOI22_X1 G1647 (
	 );
   NAND4_X1 G1646 (
	 );
   NAND3_X1 G1645 (
	 );
   NAND3_X1 G1644 (
	 );
   NAND3_X1 G1643 (
	 );
   NAND2_X1 G1642 (
	 );
   AND3_X1 G1641 (
	 );
   NAND2_X1 G1640 (
	 );
   NAND2_X1 G1639 (
	 );
   NAND4_X1 G1638 (
	 );
   NAND3_X1 G1637 (
	 );
   NAND3_X1 G1636 (
	 );
   NAND3_X1 G1635 (
	 );
   NAND2_X1 G1634 (
	 );
   NAND2_X1 G1633 (
	 );
   NAND4_X1 G1632 (
	 );
   NAND3_X1 G1631 (
	 );
   NAND3_X1 G1630 (
	 );
   NAND3_X1 G1629 (
	 );
   NAND2_X1 G1628 (
	 );
   AND3_X1 G1627 (
	 );
   NAND4_X1 G1626 (
	 );
   NAND4_X1 G1625 (
	 );
   NAND4_X1 G1624 (
	 );
   CLKBUF_X1 G1623 (
	 );
   CLKBUF_X1 G1622 (
	 );
   NAND4_X1 G1621 (
	 );
   NAND4_X1 G1620 (
	 );
   NAND4_X1 G1619 (
	 );
   NAND4_X1 G1618 (
	 );
   NOR2_X1 G1617 (
	 );
   AND2_X1 G1616 (
	 );
   NAND4_X1 G1615 (
	 );
   NAND4_X1 G1614 (
	 );
   NAND3_X1 G1613 (
	 );
   NAND3_X1 G1612 (
	 );
   NAND4_X1 G1611 (
	 );
   AOI21_X1 G1610 (
	 );
   OAI21_X1 G1609 (
	 );
   AND3_X1 G1608 (
	 );
   MUX2_X1 G1607 (
	 );
   OAI21_X1 G1606 (
	 );
   INV_X1 G1605 (
	 );
   AOI22_X1 G1604 (
	 );
   MUX2_X1 G1603 (
	 );
   CLKBUF_X1 G1602 (
	 );
   AND2_X1 G1601 (
	 );
   CLKBUF_X1 G1600 (
	 );
   CLKBUF_X1 G1599 (
	 );
   OAI21_X1 G1598 (
	 );
   NAND2_X1 G1597 (
	 );
   NOR2_X1 G1596 (
	 );
   INV_X1 G1595 (
	 );
   OAI211_X1 G1594 (
	 );
   CLKBUF_X1 G1593 (
	 );
   CLKBUF_X1 G1592 (
	 );
   CLKBUF_X1 G1591 (
	 );
   CLKBUF_X1 G1590 (
	 );
   CLKBUF_X1 G1589 (
	 );
   CLKBUF_X1 G1588 (
	 );
   CLKBUF_X1 G1587 (
	 );
   CLKBUF_X1 G1586 (
	 );
   CLKBUF_X1 G1585 (
	 );
   CLKBUF_X1 G1584 (
	 );
   CLKBUF_X1 G1583 (
	 );
   CLKBUF_X1 G1582 (
	 );
   NOR2_X1 G1581 (
	 );
   CLKBUF_X1 G1580 (
	 );
   CLKBUF_X1 G1579 (
	 );
   NOR3_X1 G1578 (
	 );
   AOI21_X1 G1577 (
	 );
   NOR3_X1 G1576 (
	 );
   INV_X1 G1575 (
	 );
   INV_X1 G1574 (
	 );
   INV_X1 G1573 (
	 );
   OAI21_X1 G1572 (
	 );
   INV_X1 G1571 (
	 );
   INV_X1 G1570 (
	 );
   NAND2_X1 G1569 (
	 );
   NAND2_X1 G1568 (
	 );
   AOI22_X1 G1567 (
	 );
   AOI22_X1 G1566 (
	 );
   OAI21_X1 G1565 (
	 );
   INV_X1 G1564 (
	 );
   NAND2_X1 G1563 (
	 );
   OAI221_X1 G1562 (
	 );
   NAND2_X1 G1561 (
	 );
   OAI21_X1 G1560 (
	 );
   INV_X1 G1559 (
	 );
   NAND2_X1 G1558 (
	 );
   CLKBUF_X1 G1557 (
	 );
   NOR2_X1 G1556 (
	 );
   NOR3_X1 G1555 (
	 );
   NOR3_X1 G1554 (
	 );
   OAI21_X1 G1553 (
	 );
   INV_X1 G1552 (
	 );
   NAND2_X1 G1551 (
	 );
   OAI22_X1 G1550 (
	 );
   CLKBUF_X1 G1549 (
	 );
   CLKBUF_X1 G1548 (
	 );
   NAND2_X1 G1547 (
	 );
   NAND2_X1 G1546 (
	 );
   NAND2_X1 G1545 (
	 );
   AOI22_X1 G1544 (
	 );
   AOI22_X1 G1543 (
	 );
   AOI22_X1 G1542 (
	 );
   NAND2_X1 G1541 (
	 );
   AOI22_X1 G1540 (
	 );
   AOI22_X1 G1539 (
	 );
   OAI21_X1 G1538 (
	 );
   NAND2_X1 G1537 (
	 );
   OAI21_X1 G1536 (
	 );
   NOR2_X1 G1535 (
	 );
   AOI21_X1 G1534 (
	 );
   INV_X1 G1533 (
	 );
   NOR2_X1 G1532 (
	 );
   NOR2_X1 G1531 (
	 );
   CLKBUF_X1 G1530 (
	 );
   CLKBUF_X1 G1529 (
	 );
   CLKBUF_X1 G1528 (
	 );
   CLKBUF_X1 G1527 (
	 );
   NOR2_X1 G1526 (
	 );
   NAND4_X1 G1525 (
	 );
   NAND2_X1 G1524 (
	 );
   AOI22_X1 G1523 (
	 );
   NAND4_X1 G1522 (
	 );
   NAND3_X1 G1521 (
	 );
   NAND3_X1 G1520 (
	 );
   NAND3_X1 G1519 (
	 );
   NAND2_X1 G1518 (
	 );
   NAND2_X1 G1517 (
	 );
   NAND2_X1 G1516 (
	 );
   NAND2_X1 G1515 (
	 );
   AOI22_X1 G1514 (
	 );
   AOI22_X1 G1513 (
	 );
   CLKBUF_X1 G1512 (
	 );
   CLKBUF_X1 G1511 (
	 );
   CLKBUF_X1 G1510 (
	 );
   MUX2_X1 G1509 (
	 );
   CLKBUF_X1 G1508 (
	 );
   MUX2_X1 G1507 (
	 );
   CLKBUF_X1 G1506 (
	 );
   OAI21_X1 G1505 (
	 );
   INV_X1 G1504 (
	 );
   OAI211_X1 G1503 (
	 );
   OAI21_X1 G1502 (
	 );
   INV_X1 G1501 (
	 );
   NAND2_X1 G1500 (
	 );
   OAI221_X1 G1499 (
	 );
   NAND2_X1 G1498 (
	 );
   CLKBUF_X1 G1497 (
	 );
   NAND2_X1 G1496 (
	 );
   AOI22_X1 G1495 (
	 );
   AOI22_X1 G1494 (
	 );
   CLKBUF_X1 G1493 (
	 );
   NAND2_X1 G1492 (
	 );
   NAND3_X1 G1491 (
	 );
   NAND2_X1 G1490 (
	 );
   INV_X1 G1489 (
	 );
   NOR2_X1 G1488 (
	 );
   AOI22_X1 G1487 (
	 );
   AOI22_X1 G1486 (
	 );
   NOR2_X1 G1485 (
	 );
   INV_X1 G1484 (
	 );
   NAND4_X1 G1483 (
	 );
   AOI22_X1 G1482 (
	 );
   NAND4_X1 G1481 (
	 );
   NAND3_X1 G1480 (
	 );
   NAND3_X1 G1479 (
	 );
   NAND3_X1 G1478 (
	 );
   NAND2_X1 G1477 (
	 );
   NAND2_X1 G1476 (
	 );
   NOR2_X1 G1475 (
	 );
   NAND2_X1 G1474 (
	 );
   NAND2_X1 G1473 (
	 );
   AOI22_X1 G1472 (
	 );
   AOI22_X1 G1471 (
	 );
   NAND2_X1 G1470 (
	 );
   NAND2_X1 G1469 (
	 );
   AOI22_X1 G1468 (
	 );
   AOI22_X1 G1467 (
	 );
   CLKBUF_X1 G1466 (
	 );
   CLKBUF_X1 G1465 (
	 );
   NOR3_X1 G1464 (
	 );
   INV_X1 G1463 (
	 );
   AOI21_X1 G1462 (
	 );
   AND3_X1 G1461 (
	 );
   CLKBUF_X1 G1460 (
	 );
   NOR4_X1 G1459 (
	 );
   INV_X1 G1458 (
	 );
   NAND2_X1 G1457 (
	 );
   INV_X1 G1456 (
	 );
   INV_X1 G1455 (
	 );
   NAND4_X1 G1454 (
	 );
   INV_X1 G1453 (
	 );
   NAND3_X1 G1452 (
	 );
   AOI22_X1 G1451 (
	 );
   NOR3_X2 G1450 (
	 );
   NAND4_X1 G1449 (
	 );
   NAND3_X1 G1448 (
	 );
   NAND3_X1 G1447 (
	 );
   NAND3_X1 G1446 (
	 );
   NAND2_X1 G1445 (
	 );
   AND3_X1 G1444 (
	 );
   NAND2_X1 G1443 (
	 );
   NAND2_X1 G1442 (
	 );
   NAND4_X1 G1441 (
	 );
   NAND3_X1 G1440 (
	 );
   NAND3_X1 G1439 (
	 );
   NAND3_X1 G1438 (
	 );
   NAND2_X1 G1437 (
	 );
   NAND2_X1 G1436 (
	 );
   NAND4_X1 G1435 (
	 );
   NAND3_X1 G1434 (
	 );
   NAND3_X1 G1433 (
	 );
   NAND3_X1 G1432 (
	 );
   NAND2_X1 G1431 (
	 );
   AND3_X1 G1430 (
	 );
   NAND4_X1 G1429 (
	 );
   BUF_X4 G1428 (
	 );
   NAND4_X1 G1427 (
	 );
   NAND4_X1 G1426 (
	 );
   BUF_X4 G1425 (
	 );
   NOR2_X1 G1424 (
	 );
   INV_X1 G1423 (
	 );
   MUX2_X1 G1422 (
	 );
   OAI21_X1 G1421 (
	 );
   INV_X1 G1420 (
	 );
   AOI22_X1 G1419 (
	 );
   NAND2_X1 G1418 (
	 );
   NAND2_X1 G1417 (
	 );
   NAND2_X1 G1416 (
	 );
   AOI22_X1 G1415 (
	 );
   AOI22_X1 G1414 (
	 );
   AOI22_X1 G1413 (
	 );
   NAND2_X1 G1412 (
	 );
   AOI22_X1 G1411 (
	 );
   AOI22_X1 G1410 (
	 );
   INV_X1 G1409 (
	 );
   MUX2_X1 G1408 (
	 );
   CLKBUF_X1 G1407 (
	 );
   OAI21_X1 G1406 (
	 );
   INV_X1 G1405 (
	 );
   NAND2_X1 G1404 (
	 );
   OAI221_X1 G1403 (
	 );
   INV_X1 G1402 (
	 );
   NAND2_X1 G1401 (
	 );
   CLKBUF_X1 G1400 (
	 );
   AND2_X1 G1399 (
	 );
   CLKBUF_X1 G1398 (
	 );
   AND2_X1 G1397 (
	 );
   AND2_X1 G1396 (
	 );
   NAND2_X1 G1395 (
	 );
   NAND2_X1 G1394 (
	 );
   NAND2_X1 G1393 (
	 );
   AOI22_X1 G1392 (
	 );
   AOI22_X1 G1391 (
	 );
   AOI22_X1 G1390 (
	 );
   NAND2_X1 G1389 (
	 );
   AOI22_X1 G1388 (
	 );
   AOI22_X1 G1387 (
	 );
   CLKBUF_X1 G1386 (
	 );
   MUX2_X1 G1385 (
	 );
   OAI21_X1 G1384 (
	 );
   INV_X1 G1383 (
	 );
   AOI22_X1 G1382 (
	 );
   CLKBUF_X1 G1381 (
	 );
   CLKBUF_X1 G1380 (
	 );
   CLKBUF_X1 G1379 (
	 );
   OAI21_X1 G1378 (
	 );
   INV_X1 G1377 (
	 );
   NAND2_X1 G1376 (
	 );
   OAI221_X1 G1375 (
	 );
   INV_X1 G1374 (
	 );
   INV_X1 G1373 (
	 );
   NAND2_X1 G1372 (
	 );
   OAI21_X1 G1371 (
	 );
   INV_X1 G1370 (
	 );
   NAND2_X1 G1369 (
	 );
   AND2_X1 G1368 (
	 );
   CLKBUF_X1 G1367 (
	 );
   AND2_X1 G1366 (
	 );
   CLKBUF_X1 G1365 (
	 );
   CLKBUF_X1 G1364 (
	 );
   CLKBUF_X1 G1363 (
	 );
   OAI21_X1 G1362 (
	 );
   INV_X1 G1361 (
	 );
   NAND2_X1 G1360 (
	 );
   CLKBUF_X1 G1359 (
	 );
   CLKBUF_X1 G1358 (
	 );
   CLKBUF_X1 G1357 (
	 );
   NOR2_X1 G1356 (
	 );
   NAND3_X1 G1355 (
	 );
   AND3_X1 G1354 (
	 );
   NAND2_X1 G1353 (
	 );
   NAND2_X1 G1352 (
	 );
   NAND2_X1 G1351 (
	 );
   AOI22_X1 G1350 (
	 );
   NAND4_X1 G1349 (
	 );
   NAND3_X1 G1348 (
	 );
   NAND3_X1 G1347 (
	 );
   NAND3_X1 G1346 (
	 );
   NAND2_X1 G1345 (
	 );
   AND3_X1 G1344 (
	 );
   NAND4_X1 G1343 (
	 );
   NAND4_X1 G1342 (
	 );
   NAND4_X1 G1341 (
	 );
   MUX2_X1 G1340 (
	 );
   OAI21_X1 G1339 (
	 );
   INV_X1 G1338 (
	 );
   NAND2_X1 G1337 (
	 );
   OAI21_X1 G1336 (
	 );
   INV_X1 G1335 (
	 );
   AOI22_X1 G1334 (
	 );
   CLKBUF_X1 G1333 (
	 );
   NAND3_X1 G1332 (
	 );
   AOI22_X1 G1331 (
	 );
   NAND4_X1 G1330 (
	 );
   NAND3_X1 G1329 (
	 );
   NAND3_X1 G1328 (
	 );
   NAND3_X1 G1327 (
	 );
   NAND2_X1 G1326 (
	 );
   AND3_X1 G1325 (
	 );
   NAND2_X1 G1324 (
	 );
   NAND2_X1 G1323 (
	 );
   NAND2_X1 G1322 (
	 );
   AND3_X1 G1321 (
	 );
   NAND4_X1 G1320 (
	 );
   NAND4_X1 G1319 (
	 );
   NAND4_X1 G1318 (
	 );
   CLKBUF_X1 G1317 (
	 );
   CLKBUF_X1 G1316 (
	 );
   OAI21_X1 G1315 (
	 );
   INV_X1 G1314 (
	 );
   NAND2_X1 G1313 (
	 );
   OAI21_X1 G1312 (
	 );
   INV_X1 G1311 (
	 );
   AOI22_X1 G1310 (
	 );
   CLKBUF_X1 G1309 (
	 );
   CLKBUF_X1 G1308 (
	 );
   CLKBUF_X1 G1307 (
	 );
   NAND4_X1 G1306 (
	 );
   NAND2_X1 G1305 (
	 );
   NAND2_X1 G1304 (
	 );
   AOI22_X1 G1303 (
	 );
   AOI22_X1 G1302 (
	 );
   NAND2_X1 G1301 (
	 );
   NAND2_X1 G1300 (
	 );
   AOI22_X1 G1299 (
	 );
   AOI22_X1 G1298 (
	 );
   NAND2_X1 G1297 (
	 );
   NOR2_X1 G1296 (
	 );
   INV_X1 G1295 (
	 );
   INV_X1 G1294 (
	 );
   AOI22_X1 G1293 (
	 );
   NAND2_X1 G1292 (
	 );
   AOI22_X1 G1291 (
	 );
   AOI22_X1 G1290 (
	 );
   CLKBUF_X1 G1289 (
	 );
   CLKBUF_X1 G1288 (
	 );
   CLKBUF_X1 G1287 (
	 );
   MUX2_X1 G1286 (
	 );
   CLKBUF_X1 G1285 (
	 );
   CLKBUF_X1 G1284 (
	 );
   CLKBUF_X1 G1283 (
	 );
   NAND2_X1 G1282 (
	 );
   AOI22_X1 G1281 (
	 );
   AOI22_X1 G1280 (
	 );
   BUF_X4 G1279 (
	 );
   CLKBUF_X1 G1278 (
	 );
   CLKBUF_X1 G1277 (
	 );
   NAND2_X1 G1276 (
	 );
   AOI22_X1 G1275 (
	 );
   AOI22_X1 G1274 (
	 );
   AND2_X1 G1273 (
	 );
   MUX2_X1 G1272 (
	 );
   OAI21_X1 G1271 (
	 );
   INV_X1 G1270 (
	 );
   NAND2_X1 G1269 (
	 );
   CLKBUF_X1 G1268 (
	 );
   MUX2_X1 G1267 (
	 );
   CLKBUF_X1 G1266 (
	 );
   CLKBUF_X1 G1265 (
	 );
   OAI21_X1 G1264 (
	 );
   INV_X1 G1263 (
	 );
   NAND2_X1 G1262 (
	 );
   OAI21_X1 G1261 (
	 );
   INV_X1 G1260 (
	 );
   AOI22_X1 G1259 (
	 );
   OAI221_X1 G1258 (
	 );
   INV_X1 G1257 (
	 );
   BUF_X4 G1256 (
	 );
   AOI22_X1 G1255 (
	 );
   INV_X1 G1254 (
	 );
   NAND2_X1 G1253 (
	 );
   CLKBUF_X1 G1252 (
	 );
   CLKBUF_X1 G1251 (
	 );
   CLKBUF_X1 G1250 (
	 );
   OAI221_X1 G1249 (
	 );
   XNOR2_X1 G1248 (
	 );
   INV_X1 G1247 (
	 );
   NAND3_X1 G1246 (
	 );
   XNOR2_X1 G1245 (
	 );
   CLKBUF_X1 G1244 (
	 );
   NAND2_X1 G1243 (
	 );
   AOI22_X1 G1242 (
	 );
   AOI22_X1 G1241 (
	 );
   BUF_X4 G1240 (
	 );
   CLKBUF_X1 G1239 (
	 );
   CLKBUF_X1 G1238 (
	 );
   CLKBUF_X1 G1237 (
	 );
   OAI21_X1 G1236 (
	 );
   INV_X1 G1235 (
	 );
   NAND2_X1 G1234 (
	 );
   OAI221_X1 G1233 (
	 );
   INV_X1 G1232 (
	 );
   INV_X1 G1231 (
	 );
   NAND2_X1 G1230 (
	 );
   CLKBUF_X1 G1229 (
	 );
   OAI221_X1 G1228 (
	 );
   NOR2_X1 G1227 (
	 );
   NAND2_X1 G1226 (
	 );
   NAND2_X1 G1225 (
	 );
   NAND4_X1 G1224 (
	 );
   NAND3_X1 G1223 (
	 );
   OAI21_X1 G1222 (
	 );
   NOR2_X1 G1221 (
	 );
   NAND2_X1 G1220 (
	 );
   INV_X1 G1219 (
	 );
   NOR2_X1 G1218 (
	 );
   NAND4_X1 G1217 (
	 );
   NAND4_X1 G1216 (
	 );
   BUF_X4 G1215 (
	 );
   NAND4_X1 G1214 (
	 );
   NAND4_X1 G1213 (
	 );
   NOR3_X1 G1212 (
	 );
   AND3_X1 G1211 (
	 );
   OAI22_X1 G1210 (
	 );
   INV_X1 G1209 (
	 );
   NAND3_X1 G1208 (
	 );
   INV_X1 G1207 (
	 );
   NAND2_X2 G1206 (
	 );
   AND2_X1 G1205 (
	 );
   INV_X1 G1204 (
	 );
   CLKBUF_X1 G1203 (
	 );
   OAI221_X1 G1202 (
	 );
   INV_X1 G1201 (
	 );
   INV_X1 G1200 (
	 );
   AOI22_X1 G1199 (
	 );
   CLKBUF_X1 G1198 (
	 );
   CLKBUF_X1 G1197 (
	 );
   NAND3_X1 G1196 (
	 );
   AOI22_X1 G1195 (
	 );
   NAND4_X1 G1194 (
	 );
   NAND3_X1 G1193 (
	 );
   NAND3_X1 G1192 (
	 );
   NAND3_X1 G1191 (
	 );
   NAND2_X1 G1190 (
	 );
   AND3_X1 G1189 (
	 );
   NAND2_X1 G1188 (
	 );
   NAND2_X1 G1187 (
	 );
   NAND4_X1 G1186 (
	 );
   NAND3_X1 G1185 (
	 );
   NAND3_X1 G1184 (
	 );
   NAND3_X1 G1183 (
	 );
   NAND2_X1 G1182 (
	 );
   NAND2_X1 G1181 (
	 );
   NAND4_X1 G1180 (
	 );
   NAND3_X1 G1179 (
	 );
   NAND3_X1 G1178 (
	 );
   NAND3_X1 G1177 (
	 );
   NAND2_X1 G1176 (
	 );
   AND3_X1 G1175 (
	 );
   NAND4_X1 G1174 (
	 );
   NAND4_X1 G1173 (
	 );
   NAND4_X1 G1172 (
	 );
   CLKBUF_X1 G1171 (
	 );
   CLKBUF_X1 G1170 (
	 );
   CLKBUF_X1 G1169 (
	 );
   MUX2_X1 G1168 (
	 );
   AOI21_X1 G1167 (
	 );
   NAND3_X1 G1166 (
	 );
   INV_X1 G1165 (
	 );
   CLKBUF_X1 G1164 (
	 );
   AOI21_X1 G1163 (
	 );
   INV_X1 G1162 (
	 );
   INV_X1 G1161 (
	 );
   CLKBUF_X1 G1160 (
	 );
   CLKBUF_X1 G1159 (
	 );
   CLKBUF_X1 G1158 (
	 );
   CLKBUF_X1 G1157 (
	 );
   CLKBUF_X1 G1156 (
	 );
   CLKBUF_X1 G1155 (
	 );
   CLKBUF_X1 G1154 (
	 );
   MUX2_X1 G1153 (
	 );
   CLKBUF_X1 G1152 (
	 );
   MUX2_X1 G1151 (
	 );
   CLKBUF_X1 G1150 (
	 );
   NOR3_X1 G1149 (
	 );
   NAND2_X1 G1148 (
	 );
   OAI21_X1 G1147 (
	 );
   INV_X1 G1146 (
	 );
   NAND2_X1 G1145 (
	 );
   OAI21_X1 G1144 (
	 );
   INV_X1 G1143 (
	 );
   AOI22_X1 G1142 (
	 );
   CLKBUF_X1 G1141 (
	 );
   OAI21_X1 G1140 (
	 );
   INV_X1 G1139 (
	 );
   NAND2_X1 G1138 (
	 );
   CLKBUF_X1 G1137 (
	 );
   AOI21_X1 G1136 (
	 );
   OAI211_X1 G1135 (
	 );
   INV_X1 G1134 (
	 );
   INV_X1 G1133 (
	 );
   OAI21_X1 G1132 (
	 );
   NOR2_X1 G1131 (
	 );
   NOR2_X1 G1130 (
	 );
   INV_X1 G1129 (
	 );
   XNOR2_X1 G1128 (
	 );
   INV_X1 G1127 (
	 );
   NAND2_X1 G1126 (
	 );
   NAND4_X1 G1125 (
	 );
   OAI21_X1 G1124 (
	 );
   OR2_X1 G1123 (
	 );
   XNOR2_X1 G1122 (
	 );
   NAND2_X1 G1121 (
	 );
   INV_X1 G1120 (
	 );
   XNOR2_X1 G1119 (
	 );
   NAND2_X1 G1118 (
	 );
   XNOR2_X1 G1117 (
	 );
   NAND3_X1 G1116 (
	 );
   AOI22_X1 G1115 (
	 );
   NOR3_X2 G1114 (
	 );
   NAND3_X1 G1113 (
	 );
   NAND4_X1 G1112 (
	 );
   NAND3_X1 G1111 (
	 );
   NAND3_X1 G1110 (
	 );
   NAND3_X1 G1109 (
	 );
   NAND2_X1 G1108 (
	 );
   BUF_X4 G1107 (
	 );
   NOR3_X1 G1106 (
	 );
   AND3_X1 G1105 (
	 );
   NAND2_X1 G1104 (
	 );
   NAND2_X1 G1103 (
	 );
   NAND4_X1 G1102 (
	 );
   NAND3_X1 G1101 (
	 );
   NAND3_X1 G1100 (
	 );
   NAND3_X1 G1099 (
	 );
   NAND2_X1 G1098 (
	 );
   NAND2_X1 G1097 (
	 );
   NAND4_X1 G1096 (
	 );
   NAND3_X1 G1095 (
	 );
   NAND3_X1 G1094 (
	 );
   BUF_X4 G1093 (
	 );
   NAND3_X1 G1092 (
	 );
   BUF_X4 G1091 (
	 );
   NAND2_X1 G1090 (
	 );
   BUF_X4 G1089 (
	 );
   AND3_X1 G1088 (
	 );
   NAND4_X1 G1087 (
	 );
   BUF_X4 G1086 (
	 );
   NAND4_X1 G1085 (
	 );
   NAND4_X1 G1084 (
	 );
   BUF_X4 G1083 (
	 );
   NOR2_X2 G1082 (
	 );
   INV_X1 G1081 (
	 );
   NOR2_X1 G1080 (
	 );
   CLKBUF_X1 G1079 (
	 );
   AND2_X1 G1078 (
	 );
   MUX2_X1 G1077 (
	 );
   OAI21_X1 G1076 (
	 );
   INV_X1 G1075 (
	 );
   AOI22_X1 G1074 (
	 );
   CLKBUF_X1 G1073 (
	 );
   CLKBUF_X1 G1072 (
	 );
   CLKBUF_X1 G1071 (
	 );
   MUX2_X1 G1070 (
	 );
   AOI21_X1 G1069 (
	 );
   AOI21_X1 G1068 (
	 );
   OAI21_X1 G1067 (
	 );
   INV_X1 G1066 (
	 );
   NOR2_X1 G1065 (
	 );
   INV_X1 G1064 (
	 );
   NAND2_X1 G1063 (
	 );
   AOI22_X1 G1062 (
	 );
   AOI22_X1 G1061 (
	 );
   CLKBUF_X1 G1060 (
	 );
   CLKBUF_X1 G1059 (
	 );
   AND2_X1 G1058 (
	 );
   MUX2_X1 G1057 (
	 );
   MUX2_X1 G1056 (
	 );
   CLKBUF_X1 G1055 (
	 );
   CLKBUF_X1 G1054 (
	 );
   CLKBUF_X1 G1053 (
	 );
   CLKBUF_X1 G1052 (
	 );
   MUX2_X1 G1051 (
	 );
   XNOR2_X1 G1050 (
	 );
   XNOR2_X1 G1049 (
	 );
   CLKBUF_X1 G1048 (
	 );
   CLKBUF_X1 G1047 (
	 );
   OAI21_X1 G1046 (
	 );
   INV_X1 G1045 (
	 );
   NAND2_X1 G1044 (
	 );
   OAI21_X1 G1043 (
	 );
   INV_X1 G1042 (
	 );
   AOI22_X1 G1041 (
	 );
   CLKBUF_X1 G1040 (
	 );
   CLKBUF_X1 G1039 (
	 );
   OAI21_X1 G1038 (
	 );
   INV_X1 G1037 (
	 );
   INV_X1 G1036 (
	 );
   NOR2_X1 G1035 (
	 );
   MUX2_X1 G1034 (
	 );
   MUX2_X1 G1033 (
	 );
   OAI21_X1 G1032 (
	 );
   INV_X1 G1031 (
	 );
   AOI22_X1 G1030 (
	 );
   CLKBUF_X1 G1029 (
	 );
   CLKBUF_X1 G1028 (
	 );
   OAI21_X1 G1027 (
	 );
   INV_X1 G1026 (
	 );
   NAND2_X1 G1025 (
	 );
   OAI21_X1 G1024 (
	 );
   INV_X1 G1023 (
	 );
   AOI22_X1 G1022 (
	 );
   CLKBUF_X1 G1021 (
	 );
   CLKBUF_X1 G1020 (
	 );
   CLKBUF_X1 G1019 (
	 );
   AND2_X1 G1018 (
	 );
   BUF_X2 G1017 (
	 );
   CLKBUF_X1 G1016 (
	 );
   AOI21_X1 G1015 (
	 );
   INV_X1 G1014 (
	 );
   CLKBUF_X1 G1013 (
	 );
   AOI21_X1 G1012 (
	 );
   INV_X1 G1011 (
	 );
   NOR2_X1 G1010 (
	 );
   BUF_X4 G1009 (
	 );
   NAND2_X2 G1008 (
	 );
   OAI21_X1 G1007 (
	 );
   BUF_X4 G1006 (
	 );
   INV_X1 G1005 (
	 );
   NAND2_X1 G1004 (
	 );
   BUF_X4 G1003 (
	 );
   BUF_X4 G1002 (
	 );
   AND2_X1 G1001 (
	 );
   NOR2_X1 G1000 (
	 );
   CLKBUF_X1 G0999 (
	 );
   CLKBUF_X1 G0998 (
	 );
   CLKBUF_X1 G0997 (
	 );
   CLKBUF_X1 G0996 (
	 );
   CLKBUF_X1 G0995 (
	 );
   CLKBUF_X1 G0994 (
	 );
   CLKBUF_X1 G0993 (
	 );
   NAND3_X1 G0992 (
	 );
   AOI22_X1 G0991 (
	 );
   AND3_X1 G0990 (
	 );
   NAND2_X1 G0989 (
	 );
   NAND2_X1 G0988 (
	 );
   NAND2_X1 G0987 (
	 );
   NAND4_X1 G0986 (
	 );
   NAND3_X1 G0985 (
	 );
   NAND3_X1 G0984 (
	 );
   NAND3_X1 G0983 (
	 );
   NAND2_X1 G0982 (
	 );
   AND3_X1 G0981 (
	 );
   NAND4_X1 G0980 (
	 );
   NAND4_X1 G0979 (
	 );
   NAND4_X1 G0978 (
	 );
   NOR2_X1 G0977 (
	 );
   CLKBUF_X1 G0976 (
	 );
   AND2_X1 G0975 (
	 );
   CLKBUF_X1 G0974 (
	 );
   NAND2_X1 G0973 (
	 );
   NAND2_X1 G0972 (
	 );
   BUF_X4 G0971 (
	 );
   NOR2_X1 G0970 (
	 );
   INV_X1 G0969 (
	 );
   NAND2_X1 G0968 (
	 );
   AOI22_X1 G0967 (
	 );
   AOI22_X1 G0966 (
	 );
   AOI22_X1 G0965 (
	 );
   BUF_X4 G0964 (
	 );
   INV_X1 G0963 (
	 );
   NAND2_X1 G0962 (
	 );
   NAND3_X1 G0961 (
	 );
   BUF_X4 G0960 (
	 );
   NOR2_X1 G0959 (
	 );
   INV_X1 G0958 (
	 );
   NAND4_X1 G0957 (
	 );
   INV_X1 G0956 (
	 );
   NAND2_X1 G0955 (
	 );
   AOI22_X1 G0954 (
	 );
   BUF_X4 G0953 (
	 );
   NOR2_X1 G0952 (
	 );
   BUF_X4 G0951 (
	 );
   NOR2_X1 G0950 (
	 );
   AOI22_X1 G0949 (
	 );
   BUF_X4 G0948 (
	 );
   NOR2_X1 G0947 (
	 );
   NOR2_X1 G0946 (
	 );
   INV_X1 G0945 (
	 );
   INV_X1 G0944 (
	 );
   CLKBUF_X1 G0943 (
	 );
   CLKBUF_X1 G0942 (
	 );
   CLKBUF_X1 G0941 (
	 );
   OAI21_X1 G0940 (
	 );
   INV_X1 G0939 (
	 );
   NAND2_X1 G0938 (
	 );
   OAI21_X1 G0937 (
	 );
   INV_X1 G0936 (
	 );
   AOI22_X1 G0935 (
	 );
   CLKBUF_X1 G0934 (
	 );
   AOI21_X1 G0933 (
	 );
   INV_X1 G0932 (
	 );
   NOR2_X1 G0931 (
	 );
   AND2_X1 G0930 (
	 );
   CLKBUF_X1 G0929 (
	 );
   AOI21_X1 G0928 (
	 );
   NAND3_X1 G0927 (
	 );
   INV_X1 G0926 (
	 );
   AND2_X2 G0925 (
	 );
   CLKBUF_X1 G0924 (
	 );
   OAI21_X1 G0923 (
	 );
   BUF_X4 G0922 (
	 );
   INV_X1 G0921 (
	 );
   NAND2_X1 G0920 (
	 );
   OAI221_X1 G0919 (
	 );
   INV_X1 G0918 (
	 );
   NAND2_X1 G0917 (
	 );
   BUF_X4 G0916 (
	 );
   BUF_X4 G0915 (
	 );
   AND2_X1 G0914 (
	 );
   NOR2_X1 G0913 (
	 );
   CLKBUF_X1 G0912 (
	 );
   CLKBUF_X1 G0911 (
	 );
   CLKBUF_X1 G0910 (
	 );
   CLKBUF_X1 G0909 (
	 );
   CLKBUF_X1 G0908 (
	 );
   CLKBUF_X1 G0907 (
	 );
   CLKBUF_X1 G0906 (
	 );
   AND2_X1 G0905 (
	 );
   AOI21_X1 G0904 (
	 );
   AOI21_X1 G0903 (
	 );
   OAI21_X1 G0902 (
	 );
   INV_X1 G0901 (
	 );
   NOR2_X1 G0900 (
	 );
   INV_X1 G0899 (
	 );
   CLKBUF_X1 G0898 (
	 );
   NAND3_X1 G0897 (
	 );
   NAND4_X1 G0896 (
	 );
   NOR3_X1 G0895 (
	 );
   NAND3_X1 G0894 (
	 );
   NAND4_X1 G0893 (
	 );
   NAND3_X1 G0892 (
	 );
   NAND3_X1 G0891 (
	 );
   OAI22_X1 G0890 (
	 );
   INV_X1 G0889 (
	 );
   INV_X1 G0888 (
	 );
   AND4_X1 G0887 (
	 );
   NOR2_X1 G0886 (
	 );
   NOR2_X1 G0885 (
	 );
   INV_X1 G0884 (
	 );
   NOR2_X1 G0883 (
	 );
   INV_X1 G0882 (
	 );
   CLKBUF_X1 G0881 (
	 );
   MUX2_X1 G0880 (
	 );
   BUF_X8 G0879 (
	 );
   NAND3_X1 G0878 (
	 );
   AND2_X1 G0877 (
	 );
   AOI21_X1 G0876 (
	 );
   INV_X1 G0875 (
	 );
   NOR2_X1 G0874 (
	 );
   NOR2_X1 G0873 (
	 );
   INV_X1 G0872 (
	 );
   AND2_X1 G0871 (
	 );
   AND2_X1 G0870 (
	 );
   NOR2_X1 G0869 (
	 );
   OAI21_X1 G0868 (
	 );
   INV_X1 G0867 (
	 );
   NAND2_X1 G0866 (
	 );
   OAI221_X1 G0865 (
	 );
   INV_X1 G0864 (
	 );
   NAND2_X1 G0863 (
	 );
   CLKBUF_X1 G0862 (
	 );
   NAND2_X1 G0861 (
	 );
   AND4_X1 G0860 (
	 );
   NAND2_X1 G0859 (
	 );
   NAND2_X1 G0858 (
	 );
   BUF_X4 G0857 (
	 );
   NOR2_X1 G0856 (
	 );
   NAND4_X1 G0855 (
	 );
   NAND3_X1 G0854 (
	 );
   NAND3_X1 G0853 (
	 );
   NAND3_X1 G0852 (
	 );
   NAND2_X1 G0851 (
	 );
   NAND2_X1 G0850 (
	 );
   NAND4_X1 G0849 (
	 );
   NAND3_X1 G0848 (
	 );
   NAND3_X1 G0847 (
	 );
   NAND3_X1 G0846 (
	 );
   NAND2_X1 G0845 (
	 );
   NAND2_X1 G0844 (
	 );
   NAND4_X1 G0843 (
	 );
   NAND3_X1 G0842 (
	 );
   NAND3_X1 G0841 (
	 );
   BUF_X4 G0840 (
	 );
   NAND3_X1 G0839 (
	 );
   BUF_X4 G0838 (
	 );
   NAND2_X1 G0837 (
	 );
   BUF_X4 G0836 (
	 );
   BUF_X4 G0835 (
	 );
   NOR3_X1 G0834 (
	 );
   AND4_X1 G0833 (
	 );
   NAND4_X1 G0832 (
	 );
   NAND4_X1 G0831 (
	 );
   BUF_X4 G0830 (
	 );
   NOR2_X2 G0829 (
	 );
   NAND3_X1 G0828 (
	 );
   NAND3_X1 G0827 (
	 );
   BUF_X4 G0826 (
	 );
   NOR3_X2 G0825 (
	 );
   INV_X1 G0824 (
	 );
   NAND2_X1 G0823 (
	 );
   INV_X1 G0822 (
	 );
   MUX2_X1 G0821 (
	 );
   CLKBUF_X1 G0820 (
	 );
   CLKBUF_X1 G0819 (
	 );
   NOR2_X1 G0818 (
	 );
   AOI21_X1 G0817 (
	 );
   MUX2_X1 G0816 (
	 );
   BUF_X8 G0815 (
	 );
   NAND2_X1 G0814 (
	 );
   NOR2_X1 G0813 (
	 );
   OAI21_X1 G0812 (
	 );
   INV_X1 G0811 (
	 );
   AOI22_X1 G0810 (
	 );
   MUX2_X1 G0809 (
	 );
   BUF_X8 G0808 (
	 );
   NAND2_X2 G0807 (
	 );
   CLKBUF_X1 G0806 (
	 );
   CLKBUF_X1 G0805 (
	 );
   OAI21_X1 G0804 (
	 );
   INV_X1 G0803 (
	 );
   NAND2_X1 G0802 (
	 );
   OAI21_X1 G0801 (
	 );
   INV_X1 G0800 (
	 );
   AOI22_X1 G0799 (
	 );
   OAI221_X1 G0798 (
	 );
   INV_X1 G0797 (
	 );
   INV_X1 G0796 (
	 );
   AOI22_X1 G0795 (
	 );
   MUX2_X1 G0794 (
	 );
   OAI21_X1 G0793 (
	 );
   INV_X1 G0792 (
	 );
   AOI22_X1 G0791 (
	 );
   CLKBUF_X1 G0790 (
	 );
   CLKBUF_X1 G0789 (
	 );
   CLKBUF_X1 G0788 (
	 );
   AOI21_X1 G0787 (
	 );
   INV_X1 G0786 (
	 );
   NAND3_X1 G0785 (
	 );
   AOI21_X1 G0784 (
	 );
   AOI21_X1 G0783 (
	 );
   OAI21_X1 G0782 (
	 );
   INV_X1 G0781 (
	 );
   NOR2_X1 G0780 (
	 );
   INV_X1 G0779 (
	 );
   INV_X1 G0778 (
	 );
   CLKBUF_X1 G0777 (
	 );
   CLKBUF_X1 G0776 (
	 );
   MUX2_X1 G0775 (
	 );
   BUF_X8 G0774 (
	 );
   NAND3_X1 G0773 (
	 );
   INV_X1 G0772 (
	 );
   OAI21_X1 G0771 (
	 );
   INV_X1 G0770 (
	 );
   AOI22_X1 G0769 (
	 );
   OAI21_X1 G0768 (
	 );
   INV_X1 G0767 (
	 );
   NAND2_X1 G0766 (
	 );
   OAI221_X1 G0765 (
	 );
   INV_X1 G0764 (
	 );
   INV_X1 G0763 (
	 );
   NAND2_X1 G0762 (
	 );
   CLKBUF_X1 G0761 (
	 );
   CLKBUF_X1 G0760 (
	 );
   CLKBUF_X1 G0759 (
	 );
   CLKBUF_X1 G0758 (
	 );
   OAI21_X1 G0757 (
	 );
   INV_X1 G0756 (
	 );
   NAND2_X1 G0755 (
	 );
   OAI221_X1 G0754 (
	 );
   INV_X1 G0753 (
	 );
   NAND2_X1 G0752 (
	 );
   CLKBUF_X1 G0751 (
	 );
   CLKBUF_X1 G0750 (
	 );
   CLKBUF_X1 G0749 (
	 );
   MUX2_X1 G0748 (
	 );
   CLKBUF_X1 G0747 (
	 );
   NOR2_X1 G0746 (
	 );
   CLKBUF_X1 G0745 (
	 );
   CLKBUF_X1 G0744 (
	 );
   NAND2_X1 G0743 (
	 );
   NAND2_X1 G0742 (
	 );
   AOI22_X1 G0741 (
	 );
   CLKBUF_X1 G0740 (
	 );
   CLKBUF_X1 G0739 (
	 );
   OAI221_X1 G0738 (
	 );
   INV_X1 G0737 (
	 );
   INV_X1 G0736 (
	 );
   AOI22_X1 G0735 (
	 );
   CLKBUF_X1 G0734 (
	 );
   CLKBUF_X1 G0733 (
	 );
   NAND2_X1 G0732 (
	 );
   AOI22_X1 G0731 (
	 );
   INV_X2 G0730 (
	 );
   AOI22_X1 G0729 (
	 );
   CLKBUF_X1 G0728 (
	 );
   MUX2_X1 G0727 (
	 );
   MUX2_X1 G0726 (
	 );
   CLKBUF_X1 G0725 (
	 );
   CLKBUF_X1 G0724 (
	 );
   NOR3_X1 G0723 (
	 );
   AOI21_X1 G0722 (
	 );
   INV_X1 G0721 (
	 );
   NAND3_X1 G0720 (
	 );
   INV_X1 G0719 (
	 );
   NOR2_X1 G0718 (
	 );
   NOR2_X1 G0717 (
	 );
   NAND2_X1 G0716 (
	 );
   INV_X1 G0715 (
	 );
   NAND4_X1 G0714 (
	 );
   INV_X1 G0713 (
	 );
   INV_X1 G0712 (
	 );
   CLKBUF_X1 G0711 (
	 );
   CLKBUF_X1 G0710 (
	 );
   AND2_X1 G0709 (
	 );
   MUX2_X1 G0708 (
	 );
   BUF_X8 G0707 (
	 );
   BUF_X8 G0706 (
	 );
   NAND2_X1 G0705 (
	 );
   CLKBUF_X1 G0704 (
	 );
   CLKBUF_X1 G0703 (
	 );
   CLKBUF_X1 G0702 (
	 );
   AOI21_X1 G0701 (
	 );
   INV_X1 G0700 (
	 );
   INV_X1 G0699 (
	 );
   BUF_X4 G0698 (
	 );
   INV_X1 G0697 (
	 );
   NAND2_X1 G0696 (
	 );
   NOR2_X2 G0695 (
	 );
   NAND3_X1 G0694 (
	 );
   INV_X1 G0693 (
	 );
   AND3_X2 G0692 (
	 );
   AND3_X1 G0691 (
	 );
   CLKBUF_X1 G0690 (
	 );
   NAND2_X1 G0689 (
	 );
   NAND2_X1 G0688 (
	 );
   NAND2_X1 G0687 (
	 );
   AOI22_X1 G0686 (
	 );
   AOI22_X1 G0685 (
	 );
   AOI22_X1 G0684 (
	 );
   NAND2_X1 G0683 (
	 );
   AOI22_X1 G0682 (
	 );
   AOI22_X1 G0681 (
	 );
   CLKBUF_X1 G0680 (
	 );
   NAND2_X1 G0679 (
	 );
   AOI22_X1 G0678 (
	 );
   AOI22_X1 G0677 (
	 );
   CLKBUF_X1 G0676 (
	 );
   NAND2_X1 G0675 (
	 );
   INV_X1 G0674 (
	 );
   NAND2_X1 G0673 (
	 );
   NAND3_X1 G0672 (
	 );
   NAND4_X1 G0671 (
	 );
   BUF_X4 G0670 (
	 );
   AND2_X2 G0669 (
	 );
   NOR3_X1 G0668 (
	 );
   NAND3_X1 G0667 (
	 );
   NAND4_X1 G0666 (
	 );
   BUF_X4 G0665 (
	 );
   NOR2_X2 G0664 (
	 );
   BUF_X4 G0663 (
	 );
   BUF_X4 G0662 (
	 );
   AND2_X1 G0661 (
	 );
   NAND3_X1 G0660 (
	 );
   BUF_X4 G0659 (
	 );
   NOR2_X2 G0658 (
	 );
   BUF_X4 G0657 (
	 );
   BUF_X4 G0656 (
	 );
   AND3_X1 G0655 (
	 );
   NAND3_X1 G0654 (
	 );
   BUF_X4 G0653 (
	 );
   NOR2_X2 G0652 (
	 );
   BUF_X4 G0651 (
	 );
   NOR3_X2 G0650 (
	 );
   OAI22_X1 G0649 (
	 );
   BUF_X4 G0648 (
	 );
   OAI211_X1 G0647 (
	 );
   INV_X1 G0646 (
	 );
   INV_X1 G0645 (
	 );
   OAI211_X2 G0644 (
	 );
   NAND3_X1 G0643 (
	 );
   AND4_X1 G0642 (
	 );
   NOR3_X2 G0641 (
	 );
   BUF_X4 G0640 (
	 );
   BUF_X4 G0639 (
	 );
   NOR2_X1 G0638 (
	 );
   NOR2_X1 G0637 (
	 );
   BUF_X4 G0636 (
	 );
   NAND4_X1 G0635 (
	 );
   NOR2_X2 G0634 (
	 );
   NOR2_X1 G0633 (
	 );
   BUF_X4 G0632 (
	 );
   NAND4_X1 G0631 (
	 );
   BUF_X4 G0630 (
	 );
   NAND4_X1 G0629 (
	 );
   INV_X1 G0628 (
	 );
   NAND4_X1 G0627 (
	 );
   INV_X1 G0626 (
	 );
   INV_X1 G0625 (
	 );
   NOR2_X2 G0624 (
	 );
   NAND2_X1 G0623 (
	 );
   AOI22_X1 G0622 (
	 );
   AOI22_X1 G0621 (
	 );
   BUF_X4 G0620 (
	 );
   CLKBUF_X1 G0619 (
	 );
   AND2_X1 G0618 (
	 );
   AND2_X1 G0617 (
	 );
   INV_X1 G0616 (
	 );
   AOI211_X1 G0615 (
	 );
   AOI21_X1 G0614 (
	 );
   OAI21_X1 G0613 (
	 );
   INV_X1 G0612 (
	 );
   NOR2_X1 G0611 (
	 );
   INV_X1 G0610 (
	 );
   INV_X1 G0609 (
	 );
   OAI21_X1 G0608 (
	 );
   INV_X1 G0607 (
	 );
   NAND2_X1 G0606 (
	 );
   OAI22_X1 G0605 (
	 );
   INV_X1 G0604 (
	 );
   INV_X1 G0603 (
	 );
   CLKBUF_X1 G0602 (
	 );
   AND2_X1 G0601 (
	 );
   AOI21_X1 G0600 (
	 );
   INV_X1 G0599 (
	 );
   NOR2_X1 G0598 (
	 );
   NOR2_X1 G0597 (
	 );
   BUF_X4 G0596 (
	 );
   NAND2_X2 G0595 (
	 );
   OAI21_X1 G0594 (
	 );
   INV_X1 G0593 (
	 );
   NAND2_X1 G0592 (
	 );
   OAI21_X1 G0591 (
	 );
   INV_X1 G0590 (
	 );
   AOI22_X1 G0589 (
	 );
   CLKBUF_X1 G0588 (
	 );
   CLKBUF_X1 G0587 (
	 );
   AND2_X1 G0586 (
	 );
   CLKBUF_X1 G0585 (
	 );
   CLKBUF_X1 G0584 (
	 );
   OAI221_X1 G0583 (
	 );
   BUF_X4 G0582 (
	 );
   INV_X1 G0581 (
	 );
   INV_X1 G0580 (
	 );
   AOI22_X1 G0579 (
	 );
   INV_X1 G0578 (
	 );
   OAI221_X1 G0577 (
	 );
   BUF_X4 G0576 (
	 );
   NAND2_X1 G0575 (
	 );
   INV_X1 G0574 (
	 );
   BUF_X4 G0573 (
	 );
   INV_X1 G0572 (
	 );
   NOR2_X2 G0571 (
	 );
   INV_X1 G0570 (
	 );
   AOI22_X1 G0569 (
	 );
   BUF_X4 G0568 (
	 );
   NOR2_X1 G0567 (
	 );
   BUF_X4 G0566 (
	 );
   AND2_X1 G0565 (
	 );
   INV_X1 G0564 (
	 );
   OAI221_X1 G0563 (
	 );
   INV_X1 G0562 (
	 );
   NAND2_X1 G0561 (
	 );
   NAND3_X1 G0560 (
	 );
   OAI21_X1 G0559 (
	 );
   OAI21_X1 G0558 (
	 );
   NOR2_X1 G0557 (
	 );
   MUX2_X1 G0556 (
	 );
   BUF_X8 G0555 (
	 );
   NAND3_X2 G0554 (
	 );
   NOR2_X1 G0553 (
	 );
   INV_X1 G0552 (
	 );
   NOR2_X1 G0551 (
	 );
   OAI21_X1 G0550 (
	 );
   BUF_X4 G0549 (
	 );
   INV_X1 G0548 (
	 );
   NAND2_X1 G0547 (
	 );
   OAI221_X1 G0546 (
	 );
   INV_X1 G0545 (
	 );
   INV_X1 G0544 (
	 );
   NAND2_X1 G0543 (
	 );
   BUF_X4 G0542 (
	 );
   BUF_X4 G0541 (
	 );
   AND2_X1 G0540 (
	 );
   NOR2_X1 G0539 (
	 );
   INV_X1 G0538 (
	 );
   CLKBUF_X1 G0537 (
	 );
   NAND2_X1 G0536 (
	 );
   INV_X1 G0535 (
	 );
   NAND2_X1 G0534 (
	 );
   AND2_X1 G0533 (
	 );
   BUF_X4 G0532 (
	 );
   CLKBUF_X1 G0531 (
	 );
   AND2_X1 G0530 (
	 );
   OAI21_X1 G0529 (
	 );
   BUF_X4 G0528 (
	 );
   INV_X1 G0527 (
	 );
   NAND2_X1 G0526 (
	 );
   OAI21_X1 G0525 (
	 );
   INV_X1 G0524 (
	 );
   AOI22_X1 G0523 (
	 );
   BUF_X4 G0522 (
	 );
   BUF_X4 G0521 (
	 );
   AND2_X1 G0520 (
	 );
   NOR2_X1 G0519 (
	 );
   INV_X1 G0518 (
	 );
   AND2_X1 G0517 (
	 );
   CLKBUF_X1 G0516 (
	 );
   CLKBUF_X1 G0515 (
	 );
   CLKBUF_X1 G0514 (
	 );
   AND2_X1 G0513 (
	 );
   CLKBUF_X1 G0512 (
	 );
   CLKBUF_X1 G0511 (
	 );
   AND2_X1 G0510 (
	 );
   BUF_X2 G0509 (
	 );
   CLKBUF_X1 G0508 (
	 );
   AOI21_X1 G0507 (
	 );
   NOR3_X1 G0506 (
	 );
   INV_X2 G0505 (
	 );
   NOR3_X1 G0504 (
	 );
   OR4_X1 G0503 (
	 );
   NOR2_X1 G0502 (
	 );
   INV_X1 G0501 (
	 );
   NAND2_X1 G0500 (
	 );
   NAND2_X1 G0499 (
	 );
   INV_X1 G0498 (
	 );
   NAND2_X1 G0497 (
	 );
   OAI21_X1 G0496 (
	 );
   BUF_X4 G0495 (
	 );
   INV_X1 G0494 (
	 );
   NAND2_X1 G0493 (
	 );
   BUF_X4 G0492 (
	 );
   BUF_X4 G0491 (
	 );
   AND2_X1 G0490 (
	 );
   NOR2_X1 G0489 (
	 );
   INV_X1 G0488 (
	 );
   MUX2_X1 G0487 (
	 );
   OAI21_X1 G0486 (
	 );
   INV_X1 G0485 (
	 );
   INV_X1 G0484 (
	 );
   NAND2_X1 G0483 (
	 );
   OAI21_X1 G0482 (
	 );
   INV_X1 G0481 (
	 );
   BUF_X4 G0480 (
	 );
   NOR2_X1 G0479 (
	 );
   INV_X1 G0478 (
	 );
   NOR2_X1 G0477 (
	 );
   NAND2_X1 G0476 (
	 );
   INV_X1 G0475 (
	 );
   NAND2_X1 G0474 (
	 );
   BUF_X4 G0473 (
	 );
   NOR2_X1 G0472 (
	 );
   INV_X1 G0471 (
	 );
   NAND4_X1 G0470 (
	 );
   INV_X1 G0469 (
	 );
   NAND2_X1 G0468 (
	 );
   AOI22_X1 G0467 (
	 );
   BUF_X4 G0466 (
	 );
   NOR2_X1 G0465 (
	 );
   BUF_X4 G0464 (
	 );
   NOR2_X1 G0463 (
	 );
   AOI22_X1 G0462 (
	 );
   BUF_X4 G0461 (
	 );
   NOR2_X1 G0460 (
	 );
   BUF_X4 G0459 (
	 );
   NOR2_X1 G0458 (
	 );
   INV_X1 G0457 (
	 );
   INV_X1 G0456 (
	 );
   NOR3_X1 G0455 (
	 );
   OR4_X1 G0454 (
	 );
   INV_X1 G0453 (
	 );
   NAND2_X1 G0452 (
	 );
   INV_X1 G0451 (
	 );
   NOR3_X1 G0450 (
	 );
   INV_X1 G0449 (
	 );
   INV_X1 G0448 (
	 );
   NAND2_X1 G0447 (
	 );
   NAND3_X1 G0446 (
	 );
   AND3_X1 G0445 (
	 );
   NAND2_X1 G0444 (
	 );
   NAND2_X1 G0443 (
	 );
   NAND4_X1 G0442 (
	 );
   NAND3_X1 G0441 (
	 );
   NAND3_X1 G0440 (
	 );
   NAND3_X1 G0439 (
	 );
   NAND2_X1 G0438 (
	 );
   NAND2_X1 G0437 (
	 );
   BUF_X4 G0436 (
	 );
   NAND4_X1 G0435 (
	 );
   NAND3_X1 G0434 (
	 );
   NAND3_X1 G0433 (
	 );
   NAND3_X1 G0432 (
	 );
   NAND2_X1 G0431 (
	 );
   AOI22_X1 G0430 (
	 );
   NAND4_X1 G0429 (
	 );
   NAND3_X1 G0428 (
	 );
   NAND3_X1 G0427 (
	 );
   NAND3_X1 G0426 (
	 );
   NAND2_X1 G0425 (
	 );
   AND3_X1 G0424 (
	 );
   NAND4_X1 G0423 (
	 );
   NAND4_X1 G0422 (
	 );
   NAND4_X1 G0421 (
	 );
   NOR2_X1 G0420 (
	 );
   NOR2_X1 G0419 (
	 );
   INV_X1 G0418 (
	 );
   CLKBUF_X1 G0417 (
	 );
   CLKBUF_X1 G0416 (
	 );
   CLKBUF_X1 G0415 (
	 );
   CLKBUF_X1 G0414 (
	 );
   CLKBUF_X1 G0413 (
	 );
   CLKBUF_X1 G0412 (
	 );
   CLKBUF_X1 G0411 (
	 );
   CLKBUF_X1 G0410 (
	 );
   CLKBUF_X1 G0409 (
	 );
   NAND3_X1 G0408 (
	 );
   AOI22_X1 G0407 (
	 );
   NOR3_X2 G0406 (
	 );
   NAND3_X1 G0405 (
	 );
   NAND4_X1 G0404 (
	 );
   NAND3_X1 G0403 (
	 );
   NAND3_X1 G0402 (
	 );
   NAND3_X1 G0401 (
	 );
   NAND2_X1 G0400 (
	 );
   AND3_X1 G0399 (
	 );
   NAND2_X1 G0398 (
	 );
   NAND2_X1 G0397 (
	 );
   NAND4_X1 G0396 (
	 );
   NAND3_X1 G0395 (
	 );
   NAND3_X1 G0394 (
	 );
   NAND3_X1 G0393 (
	 );
   NAND2_X1 G0392 (
	 );
   NAND2_X1 G0391 (
	 );
   AND3_X1 G0390 (
	 );
   NAND4_X1 G0389 (
	 );
   BUF_X4 G0388 (
	 );
   NAND4_X1 G0387 (
	 );
   NAND4_X1 G0386 (
	 );
   BUF_X4 G0385 (
	 );
   NOR2_X1 G0384 (
	 );
   INV_X1 G0383 (
	 );
   OAI21_X1 G0382 (
	 );
   BUF_X4 G0381 (
	 );
   INV_X1 G0380 (
	 );
   NAND2_X1 G0379 (
	 );
   OAI221_X1 G0378 (
	 );
   INV_X1 G0377 (
	 );
   INV_X2 G0376 (
	 );
   INV_X1 G0375 (
	 );
   INV_X1 G0374 (
	 );
   NAND2_X1 G0373 (
	 );
   BUF_X4 G0372 (
	 );
   BUF_X4 G0371 (
	 );
   BUF_X4 G0370 (
	 );
   AND2_X1 G0369 (
	 );
   INV_X1 G0368 (
	 );
   NAND2_X1 G0367 (
	 );
   CLKBUF_X1 G0366 (
	 );
   CLKBUF_X1 G0365 (
	 );
   NAND4_X1 G0364 (
	 );
   AOI22_X1 G0363 (
	 );
   BUF_X4 G0362 (
	 );
   NOR2_X1 G0361 (
	 );
   INV_X1 G0360 (
	 );
   BUF_X4 G0359 (
	 );
   NOR2_X1 G0358 (
	 );
   INV_X1 G0357 (
	 );
   NAND4_X1 G0356 (
	 );
   NAND3_X1 G0355 (
	 );
   NAND3_X1 G0354 (
	 );
   NAND3_X1 G0353 (
	 );
   NAND2_X1 G0352 (
	 );
   NAND2_X1 G0351 (
	 );
   NAND4_X1 G0350 (
	 );
   NAND3_X1 G0349 (
	 );
   NAND3_X1 G0348 (
	 );
   BUF_X4 G0347 (
	 );
   NAND3_X1 G0346 (
	 );
   BUF_X4 G0345 (
	 );
   NAND2_X1 G0344 (
	 );
   NOR2_X1 G0343 (
	 );
   INV_X1 G0342 (
	 );
   NAND2_X1 G0341 (
	 );
   BUF_X4 G0340 (
	 );
   NOR2_X1 G0339 (
	 );
   INV_X1 G0338 (
	 );
   NAND4_X1 G0337 (
	 );
   INV_X1 G0336 (
	 );
   NAND2_X1 G0335 (
	 );
   AOI22_X1 G0334 (
	 );
   BUF_X4 G0333 (
	 );
   AOI22_X1 G0332 (
	 );
   NAND2_X1 G0331 (
	 );
   BUF_X4 G0330 (
	 );
   NOR2_X1 G0329 (
	 );
   NAND3_X1 G0328 (
	 );
   NOR2_X1 G0327 (
	 );
   NOR2_X1 G0326 (
	 );
   NAND2_X1 G0325 (
	 );
   NAND2_X1 G0324 (
	 );
   AOI22_X1 G0323 (
	 );
   BUF_X4 G0322 (
	 );
   NOR2_X1 G0321 (
	 );
   BUF_X4 G0320 (
	 );
   NOR2_X1 G0319 (
	 );
   INV_X1 G0318 (
	 );
   AOI22_X1 G0317 (
	 );
   INV_X1 G0316 (
	 );
   NAND2_X1 G0315 (
	 );
   BUF_X4 G0314 (
	 );
   NOR2_X1 G0313 (
	 );
   INV_X1 G0312 (
	 );
   CLKBUF_X1 G0311 (
	 );
   CLKBUF_X1 G0310 (
	 );
   CLKBUF_X1 G0309 (
	 );
   CLKBUF_X1 G0308 (
	 );
   CLKBUF_X1 G0307 (
	 );
   NOR2_X1 G0306 (
	 );
   BUF_X4 G0305 (
	 );
   INV_X2 G0304 (
	 );
   CLKBUF_X1 G0303 (
	 );
   CLKBUF_X1 G0302 (
	 );
   CLKBUF_X1 G0301 (
	 );
   MUX2_X1 G0300 (
	 );
   BUF_X8 G0299 (
	 );
   NAND3_X1 G0298 (
	 );
   INV_X1 G0297 (
	 );
   AOI21_X1 G0296 (
	 );
   INV_X1 G0295 (
	 );
   NAND3_X1 G0294 (
	 );
   INV_X1 G0293 (
	 );
   OAI21_X1 G0292 (
	 );
   INV_X1 G0291 (
	 );
   BUF_X4 G0290 (
	 );
   INV_X2 G0289 (
	 );
   NOR2_X1 G0288 (
	 );
   AOI22_X1 G0287 (
	 );
   CLKBUF_X1 G0286 (
	 );
   NAND4_X1 G0285 (
	 );
   NAND2_X1 G0284 (
	 );
   BUF_X4 G0283 (
	 );
   NOR2_X1 G0282 (
	 );
   NAND2_X1 G0281 (
	 );
   AOI22_X1 G0280 (
	 );
   AOI22_X1 G0279 (
	 );
   NAND2_X1 G0278 (
	 );
   NAND4_X1 G0277 (
	 );
   NAND3_X1 G0276 (
	 );
   NAND3_X1 G0275 (
	 );
   BUF_X4 G0274 (
	 );
   NAND3_X1 G0273 (
	 );
   BUF_X4 G0272 (
	 );
   NAND2_X1 G0271 (
	 );
   NOR2_X1 G0270 (
	 );
   INV_X1 G0269 (
	 );
   NAND3_X1 G0268 (
	 );
   NOR2_X1 G0267 (
	 );
   NAND2_X1 G0266 (
	 );
   BUF_X4 G0265 (
	 );
   NOR2_X1 G0264 (
	 );
   INV_X1 G0263 (
	 );
   NAND2_X1 G0262 (
	 );
   AOI22_X1 G0261 (
	 );
   BUF_X4 G0260 (
	 );
   BUF_X4 G0259 (
	 );
   AOI22_X1 G0258 (
	 );
   BUF_X4 G0257 (
	 );
   AOI22_X1 G0256 (
	 );
   BUF_X4 G0255 (
	 );
   NOR2_X1 G0254 (
	 );
   INV_X1 G0253 (
	 );
   NOR2_X1 G0252 (
	 );
   NAND2_X1 G0251 (
	 );
   BUF_X4 G0250 (
	 );
   NOR2_X1 G0249 (
	 );
   INV_X1 G0248 (
	 );
   NAND4_X1 G0247 (
	 );
   INV_X1 G0246 (
	 );
   NAND2_X1 G0245 (
	 );
   AOI22_X1 G0244 (
	 );
   BUF_X4 G0243 (
	 );
   NOR2_X1 G0242 (
	 );
   NOR2_X1 G0241 (
	 );
   INV_X1 G0240 (
	 );
   AOI22_X1 G0239 (
	 );
   INV_X1 G0238 (
	 );
   NAND2_X1 G0237 (
	 );
   NOR2_X1 G0236 (
	 );
   INV_X1 G0235 (
	 );
   NAND2_X1 G0234 (
	 );
   INV_X1 G0233 (
	 );
   OAI21_X1 G0232 (
	 );
   INV_X1 G0231 (
	 );
   INV_X1 G0230 (
	 );
   INV_X1 G0229 (
	 );
   OAI21_X1 G0228 (
	 );
   BUF_X4 G0227 (
	 );
   INV_X1 G0226 (
	 );
   NAND2_X1 G0225 (
	 );
   OAI21_X1 G0224 (
	 );
   INV_X1 G0223 (
	 );
   BUF_X4 G0222 (
	 );
   INV_X1 G0221 (
	 );
   AOI22_X1 G0220 (
	 );
   BUF_X4 G0219 (
	 );
   BUF_X4 G0218 (
	 );
   AND2_X1 G0217 (
	 );
   NOR2_X1 G0216 (
	 );
   AND2_X2 G0215 (
	 );
   NAND2_X1 G0214 (
	 );
   INV_X1 G0213 (
	 );
   NOR2_X2 G0212 (
	 );
   NOR3_X1 G0211 (
	 );
   INV_X1 G0210 (
	 );
   INV_X1 G0209 (
	 );
   OAI21_X1 G0208 (
	 );
   INV_X1 G0207 (
	 );
   NAND2_X1 G0206 (
	 );
   OAI221_X1 G0205 (
	 );
   INV_X1 G0204 (
	 );
   INV_X1 G0203 (
	 );
   NAND2_X1 G0202 (
	 );
   CLKBUF_X1 G0201 (
	 );
   CLKBUF_X1 G0200 (
	 );
   CLKBUF_X1 G0199 (
	 );
   CLKBUF_X1 G0198 (
	 );
   CLKBUF_X1 G0197 (
	 );
   CLKBUF_X1 G0196 (
	 );
   CLKBUF_X1 G0195 (
	 );
   CLKBUF_X1 G0194 (
	 );
   MUX2_X1 G0193 (
	 );
   CLKBUF_X1 G0192 (
	 );
   OAI221_X1 G0191 (
	 );
   BUF_X4 G0190 (
	 );
   NAND2_X1 G0189 (
	 );
   INV_X1 G0188 (
	 );
   BUF_X4 G0187 (
	 );
   NAND2_X1 G0186 (
	 );
   INV_X1 G0185 (
	 );
   AOI22_X1 G0184 (
	 );
   BUF_X4 G0183 (
	 );
   NOR2_X1 G0182 (
	 );
   BUF_X4 G0181 (
	 );
   NOR2_X1 G0180 (
	 );
   INV_X1 G0179 (
	 );
   OAI21_X1 G0178 (
	 );
   BUF_X4 G0177 (
	 );
   INV_X1 G0176 (
	 );
   NAND2_X1 G0175 (
	 );
   OAI221_X1 G0174 (
	 );
   INV_X1 G0173 (
	 );
   INV_X2 G0172 (
	 );
   INV_X2 G0171 (
	 );
   INV_X1 G0170 (
	 );
   NAND2_X1 G0169 (
	 );
   BUF_X4 G0168 (
	 );
   BUF_X4 G0167 (
	 );
   BUF_X4 G0166 (
	 );
   AND2_X1 G0165 (
	 );
   NOR2_X1 G0164 (
	 );
   INV_X1 G0163 (
	 );
   AND2_X2 G0162 (
	 );
   NAND2_X1 G0161 (
	 );
   INV_X1 G0160 (
	 );
   NOR2_X1 G0159 (
	 );
   NOR3_X1 G0158 (
	 );
   INV_X1 G0157 (
	 );
   INV_X1 G0156 (
	 );
   CLKBUF_X1 G0155 (
	 );
   CLKBUF_X1 G0154 (
	 );
   NAND3_X1 G0153 (
	 );
   AOI22_X1 G0152 (
	 );
   NOR3_X2 G0151 (
	 );
   NAND3_X1 G0150 (
	 );
   BUF_X4 G0149 (
	 );
   NOR2_X1 G0148 (
	 );
   NAND3_X1 G0147 (
	 );
   NAND2_X1 G0146 (
	 );
   AOI22_X1 G0145 (
	 );
   AOI22_X1 G0144 (
	 );
   INV_X1 G0143 (
	 );
   NAND2_X1 G0142 (
	 );
   AND3_X1 G0141 (
	 );
   NAND2_X1 G0140 (
	 );
   BUF_X4 G0139 (
	 );
   NOR2_X1 G0138 (
	 );
   INV_X1 G0137 (
	 );
   NOR2_X1 G0136 (
	 );
   NAND2_X1 G0135 (
	 );
   NAND2_X1 G0134 (
	 );
   BUF_X4 G0133 (
	 );
   NOR2_X1 G0132 (
	 );
   INV_X1 G0131 (
	 );
   NAND4_X1 G0130 (
	 );
   NAND3_X1 G0129 (
	 );
   NAND3_X1 G0128 (
	 );
   NAND3_X1 G0127 (
	 );
   NAND2_X1 G0126 (
	 );
   NAND2_X1 G0125 (
	 );
   BUF_X4 G0124 (
	 );
   NOR2_X1 G0123 (
	 );
   INV_X1 G0122 (
	 );
   NAND4_X1 G0121 (
	 );
   NAND3_X1 G0120 (
	 );
   NAND3_X1 G0119 (
	 );
   BUF_X4 G0118 (
	 );
   NAND3_X1 G0117 (
	 );
   BUF_X4 G0116 (
	 );
   NAND2_X1 G0115 (
	 );
   BUF_X4 G0114 (
	 );
   AND3_X1 G0113 (
	 );
   NAND4_X1 G0112 (
	 );
   BUF_X4 G0111 (
	 );
   NOR2_X1 G0110 (
	 );
   INV_X1 G0109 (
	 );
   BUF_X4 G0108 (
	 );
   NAND4_X1 G0107 (
	 );
   BUF_X4 G0106 (
	 );
   NOR2_X1 G0105 (
	 );
   NAND4_X1 G0104 (
	 );
   BUF_X4 G0103 (
	 );
   NOR2_X1 G0102 (
	 );
   INV_X1 G0101 (
	 );
   BUF_X4 G0100 (
	 );
   NOR2_X1 G0099 (
	 );
   INV_X1 G0098 (
	 );
   NOR2_X1 G0097 (
	 );
   NAND4_X1 G0096 (
	 );
   INV_X1 G0095 (
	 );
   MUX2_X1 G0094 (
	 );
   NAND2_X2 G0093 (
	 );
   NOR2_X1 G0092 (
	 );
   INV_X1 G0091 (
	 );
   NOR2_X1 G0090 (
	 );
   INV_X1 G0089 (
	 );
   CLKBUF_X1 G0088 (
	 );
   CLKBUF_X1 G0087 (
	 );
   NAND3_X1 G0086 (
	 );
   AND3_X1 G0085 (
	 );
   NAND2_X1 G0084 (
	 );
   BUF_X4 G0083 (
	 );
   NOR2_X1 G0082 (
	 );
   INV_X1 G0081 (
	 );
   NAND2_X1 G0080 (
	 );
   NOR2_X1 G0079 (
	 );
   INV_X1 G0078 (
	 );
   NAND4_X1 G0077 (
	 );
   NAND3_X1 G0076 (
	 );
   NAND3_X1 G0075 (
	 );
   NAND3_X1 G0074 (
	 );
   NAND2_X1 G0073 (
	 );
   NAND2_X1 G0072 (
	 );
   BUF_X4 G0071 (
	 );
   NOR2_X1 G0070 (
	 );
   INV_X1 G0069 (
	 );
   NAND4_X1 G0068 (
	 );
   NAND3_X1 G0067 (
	 );
   NAND3_X1 G0066 (
	 );
   NAND3_X1 G0065 (
	 );
   NAND2_X1 G0064 (
	 );
   AOI22_X1 G0063 (
	 );
   NAND4_X1 G0062 (
	 );
   NAND3_X1 G0061 (
	 );
   NAND3_X1 G0060 (
	 );
   BUF_X4 G0059 (
	 );
   NAND3_X1 G0058 (
	 );
   BUF_X4 G0057 (
	 );
   NAND2_X1 G0056 (
	 );
   BUF_X4 G0055 (
	 );
   BUF_X4 G0054 (
	 );
   NOR2_X1 G0053 (
	 );
   NAND3_X1 G0052 (
	 );
   NOR2_X1 G0051 (
	 );
   NAND2_X1 G0050 (
	 );
   NOR4_X2 G0049 (
	 );
   NAND2_X1 G0048 (
	 );
   AND3_X1 G0047 (
	 );
   NAND4_X1 G0046 (
	 );
   BUF_X4 G0045 (
	 );
   NOR2_X1 G0044 (
	 );
   INV_X1 G0043 (
	 );
   BUF_X4 G0042 (
	 );
   NAND4_X1 G0041 (
	 );
   BUF_X4 G0040 (
	 );
   NOR2_X1 G0039 (
	 );
   NAND4_X1 G0038 (
	 );
   BUF_X4 G0037 (
	 );
   NOR2_X1 G0036 (
	 );
   INV_X1 G0035 (
	 );
   BUF_X4 G0034 (
	 );
   NOR2_X1 G0033 (
	 );
   INV_X1 G0032 (
	 );
   NOR2_X1 G0031 (
	 );
   NAND4_X1 G0030 (
	 );
   INV_X1 G0029 (
	 );
   CLKBUF_X1 G0028 (
	 );
   NAND2_X1 G0027 (
	 );
   AOI22_X1 G0026 (
	 );
   BUF_X4 G0025 (
	 );
   AOI22_X1 G0024 (
	 );
   NAND2_X1 G0023 (
	 );
   AOI22_X1 G0022 (
	 );
   BUF_X4 G0021 (
	 );
   NOR2_X1 G0020 (
	 );
   BUF_X4 G0019 (
	 );
   NOR2_X1 G0018 (
	 );
   AOI22_X1 G0017 (
	 );
   BUF_X4 G0016 (
	 );
   NOR2_X1 G0015 (
	 );
   INV_X1 G0014 (
	 );
   BUF_X4 G0013 (
	 );
   NOR2_X1 G0012 (
	 );
   INV_X1 G0011 (
	 );
   CLKBUF_X1 G0010 (
	 );
   CLKBUF_X1 G0009 (
	 );
   CLKBUF_X1 G0008 (
	 );
   CLKBUF_X1 G0007 (
	 );
   CLKBUF_X1 G0006 (
	 );
   CLKBUF_X1 G0005 (
	 );
   CLKBUF_X1 G0004 (
	 );
   CLKBUF_X1 G0003 (
	 );
   CLKBUF_X1 G0002 (
	 );
   OR2_X1 G0001 (
	 );
   CLKBUF_X1 G0000 (
	 );
endmodule

