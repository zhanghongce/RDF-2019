// Written by verilog_parser.py of OpenDesign Flow Database.
// Date: 2019-07-25 20:48:06
// Format: ICCAD2015 placement contest

module usb_funct (
clk,
x1418,
x1459,
x1503,
x1547,
x1598,
x1660,
x1743,
x1792,
x185142,
x1865,
x1911,
x1974,
x2027,
x2098,
x2165,
x2214,
x2278,
x2333,
x2400,
x2477,
x2531,
x2589,
x2648,
x2707,
x2767,
x2826,
x2890,
x2968,
x3022,
x3071,
x3133,
x3194,
x3249,
x3300,
x3307,
x3314,
x3320,
x3327,
x3338,
x3349,
x3360,
x3390,
x3507,
x3534,
x3558,
x3565,
x3574,
x3588,
x3599,
x3606,
x3613,
x3621,
x3632,
x3638,
x3645,
x3653,
x3683,
x3698,
x3733,
x3772,
x3828,
x3849,
x3858,
x3867,
x3889,
x3949,
x4041,
x4117,
x4209,
x4285,
x4359,
x4449,
x4520,
x4587,
x4694,
x4781,
x4851,
x4937,
x5003,
x5077,
x5143,
x5225,
x5289,
x5364,
x5427,
x5498,
x5548,
x5601,
x5647,
x5722,
x5790,
x5850,
x5901,
x5961,
x6028,
x6102,
x6157,
x6186,
x6198,
x6220,
x6241,
x6252,
x6264,
x6282,
x6303,
x6327,
x6351,
x6401,
x6445,
x6496,
x6531,
x6577,
x6599,
net_9569,
x0,
x101,
x1010,
x1029,
x1058,
x106,
x1066,
x1074,
x1095,
x1104,
x111,
x1113,
x1121,
x1129,
x1134,
x1142,
x1153,
x116,
x1161,
x1170,
x1179,
x1187,
x1192,
x1197,
x1206,
x121,
x1215,
x1223,
x1231,
x1240,
x1248,
x126,
x1262,
x1274,
x1282,
x1290,
x1298,
x1313,
x132,
x1329,
x1343,
x1357,
x1370,
x1384,
x1402,
x143,
x157,
x166,
x182,
x19,
x198,
x208,
x223,
x233,
x244,
x257,
x268,
x27,
x277,
x285,
x293,
x297,
x304,
x316,
x329,
x33,
x341,
x348,
x355,
x366,
x374,
x381,
x389,
x39,
x401,
x413,
x420,
x427,
x437,
x447,
x454,
x46,
x461,
x465,
x472,
x480,
x494,
x507,
x526,
x555,
x57,
x589,
x637,
x65,
x682,
x715,
x73,
x732,
x747,
x769,
x784,
x798,
x80,
x813,
x86,
x871,
x890,
x898,
x906,
x91,
x911,
x916,
x921,
x926,
x931,
x936,
x941,
x948,
x957,
x962,
x987
);

// Start PIs
input clk;
input x1418;
input x1459;
input x1503;
input x1547;
input x1598;
input x1660;
input x1743;
input x1792;
input x185142;
input x1865;
input x1911;
input x1974;
input x2027;
input x2098;
input x2165;
input x2214;
input x2278;
input x2333;
input x2400;
input x2477;
input x2531;
input x2589;
input x2648;
input x2707;
input x2767;
input x2826;
input x2890;
input x2968;
input x3022;
input x3071;
input x3133;
input x3194;
input x3249;
input x3300;
input x3307;
input x3314;
input x3320;
input x3327;
input x3338;
input x3349;
input x3360;
input x3390;
input x3507;
input x3534;
input x3558;
input x3565;
input x3574;
input x3588;
input x3599;
input x3606;
input x3613;
input x3621;
input x3632;
input x3638;
input x3645;
input x3653;
input x3683;
input x3698;
input x3733;
input x3772;
input x3828;
input x3849;
input x3858;
input x3867;
input x3889;
input x3949;
input x4041;
input x4117;
input x4209;
input x4285;
input x4359;
input x4449;
input x4520;
input x4587;
input x4694;
input x4781;
input x4851;
input x4937;
input x5003;
input x5077;
input x5143;
input x5225;
input x5289;
input x5364;
input x5427;
input x5498;
input x5548;
input x5601;
input x5647;
input x5722;
input x5790;
input x5850;
input x5901;
input x5961;
input x6028;
input x6102;
input x6157;
input x6186;
input x6198;
input x6220;
input x6241;
input x6252;
input x6264;
input x6282;
input x6303;
input x6327;
input x6351;
input x6401;
input x6445;
input x6496;
input x6531;
input x6577;
input x6599;

// Start POs
output net_9569;
output x0;
output x101;
output x1010;
output x1029;
output x1058;
output x106;
output x1066;
output x1074;
output x1095;
output x1104;
output x111;
output x1113;
output x1121;
output x1129;
output x1134;
output x1142;
output x1153;
output x116;
output x1161;
output x1170;
output x1179;
output x1187;
output x1192;
output x1197;
output x1206;
output x121;
output x1215;
output x1223;
output x1231;
output x1240;
output x1248;
output x126;
output x1262;
output x1274;
output x1282;
output x1290;
output x1298;
output x1313;
output x132;
output x1329;
output x1343;
output x1357;
output x1370;
output x1384;
output x1402;
output x143;
output x157;
output x166;
output x182;
output x19;
output x198;
output x208;
output x223;
output x233;
output x244;
output x257;
output x268;
output x27;
output x277;
output x285;
output x293;
output x297;
output x304;
output x316;
output x329;
output x33;
output x341;
output x348;
output x355;
output x366;
output x374;
output x381;
output x389;
output x39;
output x401;
output x413;
output x420;
output x427;
output x437;
output x447;
output x454;
output x46;
output x461;
output x465;
output x472;
output x480;
output x494;
output x507;
output x526;
output x555;
output x57;
output x589;
output x637;
output x65;
output x682;
output x715;
output x73;
output x732;
output x747;
output x769;
output x784;
output x798;
output x80;
output x813;
output x86;
output x871;
output x890;
output x898;
output x906;
output x91;
output x911;
output x916;
output x921;
output x926;
output x931;
output x936;
output x941;
output x948;
output x957;
output x962;
output x987;

// Start wires
wire clk;
wire x1418;
wire x1459;
wire x1503;
wire x1547;
wire x1598;
wire x1660;
wire x1743;
wire x1792;
wire x185142;
wire x1865;
wire x1911;
wire x1974;
wire x2027;
wire x2098;
wire x2165;
wire x2214;
wire x2278;
wire x2333;
wire x2400;
wire x2477;
wire x2531;
wire x2589;
wire x2648;
wire x2707;
wire x2767;
wire x2826;
wire x2890;
wire x2968;
wire x3022;
wire x3071;
wire x3133;
wire x3194;
wire x3249;
wire x3300;
wire x3307;
wire x3314;
wire x3320;
wire x3327;
wire x3338;
wire x3349;
wire x3360;
wire x3390;
wire x3507;
wire x3534;
wire x3558;
wire x3565;
wire x3574;
wire x3588;
wire x3599;
wire x3606;
wire x3613;
wire x3621;
wire x3632;
wire x3638;
wire x3645;
wire x3653;
wire x3683;
wire x3698;
wire x3733;
wire x3772;
wire x3828;
wire x3849;
wire x3858;
wire x3867;
wire x3889;
wire x3949;
wire x4041;
wire x4117;
wire x4209;
wire x4285;
wire x4359;
wire x4449;
wire x4520;
wire x4587;
wire x4694;
wire x4781;
wire x4851;
wire x4937;
wire x5003;
wire x5077;
wire x5143;
wire x5225;
wire x5289;
wire x5364;
wire x5427;
wire x5498;
wire x5548;
wire x5601;
wire x5647;
wire x5722;
wire x5790;
wire x5850;
wire x5901;
wire x5961;
wire x6028;
wire x6102;
wire x6157;
wire x6186;
wire x6198;
wire x6220;
wire x6241;
wire x6252;
wire x6264;
wire x6282;
wire x6303;
wire x6327;
wire x6351;
wire x6401;
wire x6445;
wire x6496;
wire x6531;
wire x6577;
wire x6599;
wire net_9569;
wire x0;
wire x101;
wire x1010;
wire x1029;
wire x1058;
wire x106;
wire x1066;
wire x1074;
wire x1095;
wire x1104;
wire x111;
wire x1113;
wire x1121;
wire x1129;
wire x1134;
wire x1142;
wire x1153;
wire x116;
wire x1161;
wire x1170;
wire x1179;
wire x1187;
wire x1192;
wire x1197;
wire x1206;
wire x121;
wire x1215;
wire x1223;
wire x1231;
wire x1240;
wire x1248;
wire x126;
wire x1262;
wire x1274;
wire x1282;
wire x1290;
wire x1298;
wire x1313;
wire x132;
wire x1329;
wire x1343;
wire x1357;
wire x1370;
wire x1384;
wire x1402;
wire x143;
wire x157;
wire x166;
wire x182;
wire x19;
wire x198;
wire x208;
wire x223;
wire x233;
wire x244;
wire x257;
wire x268;
wire x27;
wire x277;
wire x285;
wire x293;
wire x297;
wire x304;
wire x316;
wire x329;
wire x33;
wire x341;
wire x348;
wire x355;
wire x366;
wire x374;
wire x381;
wire x389;
wire x39;
wire x401;
wire x413;
wire x420;
wire x427;
wire x437;
wire x447;
wire x454;
wire x46;
wire x461;
wire x465;
wire x472;
wire x480;
wire x494;
wire x507;
wire x526;
wire x555;
wire x57;
wire x589;
wire x637;
wire x65;
wire x682;
wire x715;
wire x73;
wire x732;
wire x747;
wire x769;
wire x784;
wire x798;
wire x80;
wire x813;
wire x86;
wire x871;
wire x890;
wire x898;
wire x906;
wire x91;
wire x911;
wire x916;
wire x921;
wire x926;
wire x931;
wire x936;
wire x941;
wire x948;
wire x957;
wire x962;
wire x987;
wire _net_10025;
wire _net_10026;
wire _net_10027;
wire _net_10028;
wire _net_10029;
wire _net_10030;
wire _net_10031;
wire _net_10032;
wire _net_10033;
wire _net_10037;
wire _net_10040;
wire _net_10041;
wire _net_10042;
wire _net_10043;
wire _net_10048;
wire _net_10049;
wire _net_10054;
wire _net_10055;
wire _net_10056;
wire _net_10057;
wire _net_10061;
wire _net_10062;
wire _net_10090;
wire _net_10091;
wire _net_10092;
wire _net_10094;
wire _net_10095;
wire _net_10096;
wire _net_10097;
wire _net_10098;
wire _net_10099;
wire _net_10100;
wire _net_10101;
wire _net_10102;
wire _net_10103;
wire _net_10104;
wire _net_10105;
wire _net_10106;
wire _net_10107;
wire _net_10108;
wire _net_10109;
wire _net_10110;
wire _net_10111;
wire _net_10112;
wire _net_10113;
wire _net_10114;
wire _net_10115;
wire _net_10116;
wire _net_10117;
wire _net_10118;
wire _net_10119;
wire _net_10120;
wire _net_10121;
wire _net_10122;
wire _net_10123;
wire _net_10124;
wire _net_10125;
wire _net_10126;
wire _net_10127;
wire _net_10128;
wire _net_10129;
wire _net_10130;
wire _net_10131;
wire _net_10136;
wire _net_10137;
wire _net_10138;
wire _net_10139;
wire _net_10140;
wire _net_10141;
wire _net_10142;
wire _net_10143;
wire _net_10144;
wire _net_10145;
wire _net_10146;
wire _net_10147;
wire _net_10148;
wire _net_10149;
wire _net_10150;
wire _net_10151;
wire _net_10152;
wire _net_10153;
wire _net_10154;
wire _net_10155;
wire _net_10156;
wire _net_10157;
wire _net_10158;
wire _net_10159;
wire _net_10160;
wire _net_10161;
wire _net_10162;
wire _net_10163;
wire _net_10164;
wire _net_10165;
wire _net_10166;
wire _net_10167;
wire _net_10168;
wire _net_10171;
wire _net_10172;
wire _net_10173;
wire _net_10174;
wire _net_10196;
wire _net_10197;
wire _net_10200;
wire _net_10201;
wire _net_10202;
wire _net_10203;
wire _net_10204;
wire _net_10205;
wire _net_10206;
wire _net_10207;
wire _net_10208;
wire _net_10209;
wire _net_10210;
wire _net_10211;
wire _net_10212;
wire _net_10213;
wire _net_10214;
wire _net_10215;
wire _net_10216;
wire _net_10217;
wire _net_10218;
wire _net_10219;
wire _net_10220;
wire _net_10221;
wire _net_10222;
wire _net_10223;
wire _net_10224;
wire _net_10225;
wire _net_10226;
wire _net_10227;
wire _net_10228;
wire _net_10229;
wire _net_10230;
wire _net_10231;
wire _net_10232;
wire _net_10233;
wire _net_10234;
wire _net_10235;
wire _net_10236;
wire _net_10241;
wire _net_10242;
wire _net_10243;
wire _net_10244;
wire _net_10245;
wire _net_10246;
wire _net_10247;
wire _net_10248;
wire _net_10249;
wire _net_10250;
wire _net_10251;
wire _net_10252;
wire _net_10253;
wire _net_10254;
wire _net_10255;
wire _net_10256;
wire _net_10257;
wire _net_10258;
wire _net_10259;
wire _net_10260;
wire _net_10261;
wire _net_10262;
wire _net_10263;
wire _net_10264;
wire _net_10265;
wire _net_10266;
wire _net_10267;
wire _net_10268;
wire _net_10269;
wire _net_10270;
wire _net_10271;
wire _net_10272;
wire _net_10273;
wire _net_10276;
wire _net_10277;
wire _net_10278;
wire _net_10279;
wire _net_10301;
wire _net_10302;
wire _net_10305;
wire _net_10306;
wire _net_10307;
wire _net_10308;
wire _net_10309;
wire _net_10310;
wire _net_10311;
wire _net_10312;
wire _net_10313;
wire _net_10314;
wire _net_10315;
wire _net_10316;
wire _net_10317;
wire _net_10318;
wire _net_10319;
wire _net_10320;
wire _net_10321;
wire _net_10322;
wire _net_10323;
wire _net_10324;
wire _net_10325;
wire _net_10326;
wire _net_10327;
wire _net_10328;
wire _net_10329;
wire _net_10330;
wire _net_10331;
wire _net_10332;
wire _net_10333;
wire _net_10334;
wire _net_10335;
wire _net_10336;
wire _net_10337;
wire _net_10338;
wire _net_10339;
wire _net_10340;
wire _net_10341;
wire _net_10346;
wire _net_10347;
wire _net_10348;
wire _net_10349;
wire _net_10350;
wire _net_10351;
wire _net_10352;
wire _net_10353;
wire _net_10354;
wire _net_10355;
wire _net_10356;
wire _net_10357;
wire _net_10358;
wire _net_10359;
wire _net_10360;
wire _net_10361;
wire _net_10362;
wire _net_10363;
wire _net_10364;
wire _net_10365;
wire _net_10366;
wire _net_10367;
wire _net_10368;
wire _net_10369;
wire _net_10370;
wire _net_10371;
wire _net_10372;
wire _net_10373;
wire _net_10374;
wire _net_10375;
wire _net_10376;
wire _net_10377;
wire _net_10378;
wire _net_10381;
wire _net_10382;
wire _net_10383;
wire _net_10384;
wire _net_10406;
wire _net_10407;
wire _net_10410;
wire _net_10411;
wire _net_10412;
wire _net_10413;
wire _net_10414;
wire _net_10415;
wire _net_10416;
wire _net_10417;
wire _net_10418;
wire _net_10419;
wire _net_10420;
wire _net_10421;
wire _net_10422;
wire _net_10423;
wire _net_10424;
wire _net_10425;
wire _net_10426;
wire _net_10427;
wire _net_10428;
wire _net_10429;
wire _net_10430;
wire _net_10431;
wire _net_10432;
wire _net_10433;
wire _net_10434;
wire _net_10435;
wire _net_10436;
wire _net_10437;
wire _net_10438;
wire _net_10439;
wire _net_10440;
wire _net_10441;
wire _net_10442;
wire _net_10443;
wire _net_10444;
wire _net_10445;
wire _net_10446;
wire _net_10451;
wire _net_10452;
wire _net_10453;
wire _net_10454;
wire _net_10455;
wire _net_10456;
wire _net_10457;
wire _net_10458;
wire _net_10459;
wire _net_10460;
wire _net_10461;
wire _net_10462;
wire _net_10463;
wire _net_10464;
wire _net_10465;
wire _net_10466;
wire _net_10467;
wire _net_10468;
wire _net_10469;
wire _net_10470;
wire _net_10471;
wire _net_10472;
wire _net_10473;
wire _net_10474;
wire _net_10475;
wire _net_10476;
wire _net_10477;
wire _net_10478;
wire _net_10479;
wire _net_10480;
wire _net_10481;
wire _net_10482;
wire _net_10483;
wire _net_10486;
wire _net_10487;
wire _net_10488;
wire _net_10489;
wire _net_10511;
wire _net_10512;
wire _net_10515;
wire _net_10528;
wire _net_10529;
wire _net_10531;
wire _net_10534;
wire _net_10535;
wire _net_10538;
wire _net_10543;
wire _net_117;
wire _net_118;
wire _net_119;
wire _net_120;
wire _net_121;
wire _net_122;
wire _net_123;
wire _net_124;
wire _net_125;
wire _net_126;
wire _net_127;
wire _net_128;
wire _net_129;
wire _net_130;
wire _net_131;
wire _net_132;
wire _net_133;
wire _net_151;
wire _net_152;
wire _net_153;
wire _net_154;
wire _net_155;
wire _net_156;
wire _net_157;
wire _net_158;
wire _net_159;
wire _net_160;
wire _net_161;
wire _net_162;
wire _net_163;
wire _net_164;
wire _net_165;
wire _net_166;
wire _net_167;
wire _net_168;
wire _net_169;
wire _net_170;
wire _net_171;
wire _net_172;
wire _net_173;
wire _net_174;
wire _net_175;
wire _net_176;
wire _net_177;
wire _net_178;
wire _net_179;
wire _net_180;
wire _net_181;
wire _net_182;
wire _net_183;
wire _net_184;
wire _net_185;
wire _net_187;
wire _net_188;
wire _net_189;
wire _net_190;
wire _net_191;
wire _net_193;
wire _net_198;
wire _net_199;
wire _net_200;
wire _net_201;
wire _net_202;
wire _net_231;
wire _net_232;
wire _net_233;
wire _net_234;
wire _net_254;
wire _net_255;
wire _net_259;
wire _net_261;
wire _net_265;
wire _net_266;
wire _net_267;
wire _net_268;
wire _net_269;
wire _net_270;
wire _net_271;
wire _net_272;
wire _net_273;
wire _net_274;
wire _net_275;
wire _net_276;
wire _net_277;
wire _net_278;
wire _net_280;
wire _net_314;
wire _net_8817;
wire _net_8819;
wire _net_8821;
wire _net_8823;
wire _net_8824;
wire _net_8825;
wire _net_8826;
wire _net_8828;
wire _net_8829;
wire _net_8830;
wire _net_8831;
wire _net_8833;
wire _net_8834;
wire _net_8839;
wire _net_8840;
wire _net_8841;
wire _net_8842;
wire _net_8843;
wire _net_8844;
wire _net_8845;
wire _net_8846;
wire _net_8847;
wire _net_8869;
wire _net_8955;
wire _net_9040;
wire _net_9062;
wire _net_9117;
wire _net_9118;
wire _net_9160;
wire _net_9161;
wire _net_9164;
wire _net_9165;
wire _net_9166;
wire _net_9167;
wire _net_9168;
wire _net_9169;
wire _net_9171;
wire _net_9172;
wire _net_9173;
wire _net_9176;
wire _net_9177;
wire _net_9178;
wire _net_9183;
wire _net_9185;
wire _net_9186;
wire _net_9187;
wire _net_9188;
wire _net_9189;
wire _net_9190;
wire _net_9191;
wire _net_9192;
wire _net_9193;
wire _net_9194;
wire _net_9195;
wire _net_9196;
wire _net_9201;
wire _net_9202;
wire _net_9203;
wire _net_9204;
wire _net_9207;
wire _net_9209;
wire _net_9211;
wire _net_9213;
wire _net_9214;
wire _net_9215;
wire _net_9217;
wire _net_9232;
wire _net_9235;
wire _net_9236;
wire _net_9237;
wire _net_9238;
wire _net_9239;
wire _net_9240;
wire _net_9241;
wire _net_9242;
wire _net_9243;
wire _net_9244;
wire _net_9245;
wire _net_9246;
wire _net_9247;
wire _net_9248;
wire _net_9249;
wire _net_9250;
wire _net_9258;
wire _net_9266;
wire _net_9267;
wire _net_9268;
wire _net_9272;
wire _net_9290;
wire _net_9291;
wire _net_9292;
wire _net_9293;
wire _net_9294;
wire _net_9295;
wire _net_9296;
wire _net_9297;
wire _net_9298;
wire _net_9299;
wire _net_9300;
wire _net_9301;
wire _net_9302;
wire _net_9309;
wire _net_9311;
wire _net_9312;
wire _net_9313;
wire _net_9314;
wire _net_9315;
wire _net_9316;
wire _net_9317;
wire _net_9318;
wire _net_9319;
wire _net_9320;
wire _net_9321;
wire _net_9322;
wire _net_9323;
wire _net_9324;
wire _net_9325;
wire _net_9326;
wire _net_9343;
wire _net_9344;
wire _net_9345;
wire _net_9346;
wire _net_9351;
wire _net_9352;
wire _net_9353;
wire _net_9354;
wire _net_9355;
wire _net_9356;
wire _net_9362;
wire _net_9363;
wire _net_9370;
wire _net_9371;
wire _net_9372;
wire _net_9373;
wire _net_9374;
wire _net_9375;
wire _net_9376;
wire _net_9377;
wire _net_9378;
wire _net_9380;
wire _net_9381;
wire _net_9382;
wire _net_9383;
wire _net_9384;
wire _net_9385;
wire _net_9386;
wire _net_9388;
wire _net_9389;
wire _net_9390;
wire _net_9391;
wire _net_9392;
wire _net_9393;
wire _net_9394;
wire _net_9395;
wire _net_9396;
wire _net_9397;
wire _net_9398;
wire _net_9399;
wire _net_9400;
wire _net_9401;
wire _net_9402;
wire _net_9403;
wire _net_9404;
wire _net_9405;
wire _net_9406;
wire _net_9407;
wire _net_9408;
wire _net_9409;
wire _net_9410;
wire _net_9411;
wire _net_9412;
wire _net_9413;
wire _net_9414;
wire _net_9415;
wire _net_9416;
wire _net_9417;
wire _net_9418;
wire _net_9419;
wire _net_9420;
wire _net_9421;
wire _net_9422;
wire _net_9423;
wire _net_9424;
wire _net_9427;
wire _net_9428;
wire _net_9429;
wire _net_9434;
wire _net_9437;
wire _net_9502;
wire _net_9503;
wire _net_9512;
wire _net_9514;
wire _net_9515;
wire _net_9516;
wire _net_9517;
wire _net_9518;
wire _net_9519;
wire _net_9520;
wire _net_9521;
wire _net_9530;
wire _net_9532;
wire _net_9536;
wire _net_9537;
wire _net_9541;
wire _net_9546;
wire _net_9547;
wire _net_9548;
wire _net_9550;
wire _net_9551;
wire _net_9552;
wire _net_9553;
wire _net_9554;
wire _net_9555;
wire _net_9556;
wire _net_9557;
wire _net_9558;
wire _net_9561;
wire _net_9562;
wire _net_9563;
wire _net_9564;
wire _net_9565;
wire _net_9566;
wire _net_9567;
wire _net_9572;
wire _net_9573;
wire _net_9580;
wire _net_9581;
wire _net_9588;
wire _net_9589;
wire _net_9590;
wire _net_9591;
wire _net_9600;
wire _net_9601;
wire _net_9602;
wire _net_9603;
wire _net_9606;
wire _net_9608;
wire _net_9609;
wire _net_9611;
wire _net_9627;
wire _net_9628;
wire _net_9629;
wire _net_9630;
wire _net_9633;
wire _net_9635;
wire _net_9636;
wire _net_9637;
wire _net_9638;
wire _net_9639;
wire _net_9640;
wire _net_9641;
wire _net_9642;
wire _net_9643;
wire _net_9644;
wire _net_9645;
wire _net_9646;
wire _net_9649;
wire _net_9658;
wire _net_9660;
wire _net_9661;
wire _net_9728;
wire _net_9729;
wire _net_9730;
wire _net_9731;
wire _net_9732;
wire _net_9733;
wire _net_9734;
wire _net_9735;
wire _net_9736;
wire _net_9740;
wire _net_9743;
wire _net_9744;
wire _net_9745;
wire _net_9746;
wire _net_9751;
wire _net_9752;
wire _net_9827;
wire _net_9828;
wire _net_9829;
wire _net_9830;
wire _net_9831;
wire _net_9832;
wire _net_9833;
wire _net_9834;
wire _net_9835;
wire _net_9839;
wire _net_9842;
wire _net_9843;
wire _net_9844;
wire _net_9845;
wire _net_9850;
wire _net_9851;
wire _net_9926;
wire _net_9927;
wire _net_9928;
wire _net_9929;
wire _net_9930;
wire _net_9931;
wire _net_9932;
wire _net_9933;
wire _net_9934;
wire _net_9938;
wire _net_9941;
wire _net_9942;
wire _net_9943;
wire _net_9944;
wire _net_9949;
wire _net_9950;
wire _net_9957;
wire _net_9958;
wire n10001;
wire n10002;
wire n10003;
wire n10004;
wire n10005;
wire n10007;
wire n10008;
wire n10009;
wire n10010;
wire n10011;
wire n10012;
wire n10013;
wire n10014;
wire n10016;
wire n10018;
wire n10019;
wire n1002;
wire n10020;
wire n10022;
wire n10024;
wire n10025;
wire n10027;
wire n10029;
wire n10030;
wire n10031;
wire n10033;
wire n10034;
wire n10035;
wire n10037;
wire n10039;
wire n10042;
wire n10043;
wire n10044;
wire n10045;
wire n10046;
wire n10047;
wire n10048;
wire n10049;
wire n10051;
wire n10055;
wire n10056;
wire n10057;
wire n10058;
wire n10059;
wire n10060;
wire n10061;
wire n10062;
wire n10063;
wire n10064;
wire n10065;
wire n10066;
wire n10067;
wire n10068;
wire n10069;
wire n1007;
wire n10071;
wire n10072;
wire n10073;
wire n10075;
wire n10076;
wire n10077;
wire n10079;
wire n10080;
wire n10081;
wire n10083;
wire n10084;
wire n10086;
wire n10087;
wire n10088;
wire n10089;
wire n10090;
wire n10091;
wire n10092;
wire n10093;
wire n10094;
wire n10095;
wire n10096;
wire n10097;
wire n10098;
wire n10099;
wire n10100;
wire n10101;
wire n10103;
wire n10104;
wire n10106;
wire n10107;
wire n10108;
wire n10109;
wire n10110;
wire n10111;
wire n10112;
wire n10113;
wire n10114;
wire n10115;
wire n10116;
wire n10117;
wire n10118;
wire n10119;
wire n1012;
wire n10120;
wire n10121;
wire n10122;
wire n10124;
wire n10126;
wire n10127;
wire n10128;
wire n10129;
wire n10130;
wire n10131;
wire n10132;
wire n10133;
wire n10134;
wire n10135;
wire n10137;
wire n10138;
wire n10140;
wire n10141;
wire n10142;
wire n10143;
wire n10144;
wire n10145;
wire n10146;
wire n10147;
wire n10148;
wire n10150;
wire n10151;
wire n10152;
wire n10153;
wire n10154;
wire n10155;
wire n10156;
wire n10157;
wire n10158;
wire n10159;
wire n10160;
wire n10161;
wire n10162;
wire n10163;
wire n10164;
wire n10165;
wire n10166;
wire n10167;
wire n10168;
wire n10169;
wire n1017;
wire n10170;
wire n10171;
wire n10172;
wire n10173;
wire n10174;
wire n10175;
wire n10176;
wire n10177;
wire n10178;
wire n10179;
wire n10180;
wire n10181;
wire n10182;
wire n10183;
wire n10185;
wire n10186;
wire n10187;
wire n10190;
wire n10191;
wire n10193;
wire n10194;
wire n10195;
wire n10196;
wire n10197;
wire n10198;
wire n10199;
wire n10201;
wire n10203;
wire n10204;
wire n10205;
wire n10207;
wire n10209;
wire n10210;
wire n10211;
wire n10213;
wire n10214;
wire n10216;
wire n10217;
wire n10219;
wire n1022;
wire n10220;
wire n10223;
wire n10224;
wire n10225;
wire n10226;
wire n10227;
wire n10229;
wire n10230;
wire n10231;
wire n10232;
wire n10233;
wire n10234;
wire n10237;
wire n10238;
wire n10239;
wire n10240;
wire n10241;
wire n10242;
wire n10243;
wire n10244;
wire n10245;
wire n10246;
wire n10247;
wire n10248;
wire n10249;
wire n10250;
wire n10251;
wire n10252;
wire n10253;
wire n10254;
wire n10255;
wire n10256;
wire n10257;
wire n10258;
wire n10259;
wire n10260;
wire n10261;
wire n10262;
wire n10263;
wire n10264;
wire n10265;
wire n10266;
wire n10267;
wire n10268;
wire n10269;
wire n1027;
wire n10271;
wire n10272;
wire n10275;
wire n10278;
wire n10279;
wire n10281;
wire n10282;
wire n10284;
wire n10285;
wire n10286;
wire n10288;
wire n10289;
wire n10290;
wire n10292;
wire n10293;
wire n10294;
wire n10295;
wire n10296;
wire n10297;
wire n10298;
wire n10299;
wire n10300;
wire n10301;
wire n10302;
wire n10303;
wire n10304;
wire n10305;
wire n10306;
wire n10307;
wire n10308;
wire n10309;
wire n10310;
wire n10311;
wire n10312;
wire n10313;
wire n10314;
wire n10315;
wire n10317;
wire n10318;
wire n10319;
wire n1032;
wire n10321;
wire n10322;
wire n10323;
wire n10325;
wire n10326;
wire n10327;
wire n10328;
wire n10329;
wire n10330;
wire n10331;
wire n10332;
wire n10334;
wire n10336;
wire n10338;
wire n10339;
wire n10340;
wire n10341;
wire n10342;
wire n10343;
wire n10344;
wire n10345;
wire n10346;
wire n10347;
wire n10348;
wire n10349;
wire n10350;
wire n10352;
wire n10353;
wire n10355;
wire n10356;
wire n10357;
wire n10358;
wire n10359;
wire n10360;
wire n10361;
wire n10362;
wire n10364;
wire n10365;
wire n10366;
wire n10367;
wire n10368;
wire n10369;
wire n1037;
wire n10370;
wire n10371;
wire n10372;
wire n10373;
wire n10375;
wire n10376;
wire n10377;
wire n10378;
wire n10379;
wire n10380;
wire n10381;
wire n10382;
wire n10383;
wire n10384;
wire n10385;
wire n10386;
wire n10387;
wire n10388;
wire n10389;
wire n10390;
wire n10391;
wire n10392;
wire n10393;
wire n10394;
wire n10395;
wire n10396;
wire n10397;
wire n10398;
wire n10399;
wire n10400;
wire n10401;
wire n10403;
wire n10404;
wire n10405;
wire n10406;
wire n10408;
wire n10409;
wire n10411;
wire n10412;
wire n10414;
wire n10415;
wire n10417;
wire n10418;
wire n10419;
wire n1042;
wire n10421;
wire n10422;
wire n10423;
wire n10424;
wire n10425;
wire n10426;
wire n10427;
wire n10428;
wire n10430;
wire n10431;
wire n10432;
wire n10433;
wire n10434;
wire n10435;
wire n10437;
wire n10438;
wire n10441;
wire n10443;
wire n10446;
wire n10447;
wire n10449;
wire n10450;
wire n10452;
wire n10453;
wire n10454;
wire n10456;
wire n10458;
wire n10459;
wire n10460;
wire n10462;
wire n10463;
wire n10464;
wire n10466;
wire n10467;
wire n10468;
wire n10469;
wire n1047;
wire n10470;
wire n10471;
wire n10472;
wire n10473;
wire n10474;
wire n10475;
wire n10476;
wire n10477;
wire n10478;
wire n10479;
wire n10480;
wire n10481;
wire n10483;
wire n10484;
wire n10485;
wire n10486;
wire n10488;
wire n10489;
wire n10490;
wire n10492;
wire n10493;
wire n10494;
wire n10495;
wire n10496;
wire n10497;
wire n10498;
wire n10499;
wire n10500;
wire n10501;
wire n10503;
wire n10504;
wire n10506;
wire n10507;
wire n10509;
wire n10510;
wire n10511;
wire n10513;
wire n10514;
wire n10516;
wire n10517;
wire n10518;
wire n1052;
wire n10520;
wire n10522;
wire n10523;
wire n10524;
wire n10525;
wire n10526;
wire n10528;
wire n10529;
wire n10530;
wire n10531;
wire n10532;
wire n10533;
wire n10534;
wire n10535;
wire n10536;
wire n10537;
wire n10538;
wire n10539;
wire n10540;
wire n10541;
wire n10542;
wire n10543;
wire n10544;
wire n10545;
wire n10546;
wire n10547;
wire n10549;
wire n10551;
wire n10552;
wire n10554;
wire n10556;
wire n10557;
wire n10559;
wire n10560;
wire n10561;
wire n10562;
wire n10563;
wire n10564;
wire n10565;
wire n10566;
wire n10567;
wire n10568;
wire n1057;
wire n10570;
wire n10571;
wire n10572;
wire n10573;
wire n10574;
wire n10575;
wire n10576;
wire n10577;
wire n10579;
wire n10580;
wire n10581;
wire n10583;
wire n10584;
wire n10586;
wire n10588;
wire n10589;
wire n10592;
wire n10593;
wire n10595;
wire n10596;
wire n10597;
wire n10598;
wire n10599;
wire n10600;
wire n10601;
wire n10603;
wire n10604;
wire n10605;
wire n10606;
wire n10607;
wire n10608;
wire n10609;
wire n10610;
wire n10611;
wire n10612;
wire n10613;
wire n10614;
wire n10615;
wire n10616;
wire n10617;
wire n1062;
wire n10620;
wire n10621;
wire n10622;
wire n10624;
wire n10625;
wire n10626;
wire n10628;
wire n10629;
wire n10630;
wire n10632;
wire n10634;
wire n10635;
wire n10636;
wire n10637;
wire n10638;
wire n10639;
wire n10640;
wire n10641;
wire n10642;
wire n10643;
wire n10644;
wire n10645;
wire n10646;
wire n10647;
wire n10648;
wire n10649;
wire n10650;
wire n10651;
wire n10652;
wire n10653;
wire n10654;
wire n10655;
wire n10656;
wire n10657;
wire n10658;
wire n10659;
wire n10660;
wire n10661;
wire n10662;
wire n10663;
wire n10664;
wire n10665;
wire n10666;
wire n10668;
wire n10669;
wire n1067;
wire n10670;
wire n10671;
wire n10672;
wire n10673;
wire n10674;
wire n10676;
wire n10677;
wire n10678;
wire n10679;
wire n10680;
wire n10681;
wire n10682;
wire n10684;
wire n10685;
wire n10686;
wire n10687;
wire n10691;
wire n10693;
wire n10694;
wire n10695;
wire n10696;
wire n10697;
wire n10698;
wire n10699;
wire n10700;
wire n10701;
wire n10702;
wire n10703;
wire n10704;
wire n10705;
wire n10706;
wire n10708;
wire n10709;
wire n10711;
wire n10713;
wire n10715;
wire n10717;
wire n10718;
wire n10719;
wire n1072;
wire n10720;
wire n10721;
wire n10722;
wire n10724;
wire n10725;
wire n10727;
wire n10728;
wire n10729;
wire n10730;
wire n10731;
wire n10732;
wire n10734;
wire n10735;
wire n10736;
wire n10738;
wire n10741;
wire n10744;
wire n10748;
wire n10749;
wire n10751;
wire n10752;
wire n10753;
wire n10755;
wire n10756;
wire n10758;
wire n10760;
wire n10762;
wire n10763;
wire n10764;
wire n10765;
wire n10766;
wire n10768;
wire n10769;
wire n1077;
wire n10770;
wire n10772;
wire n10773;
wire n10775;
wire n10776;
wire n10777;
wire n10779;
wire n10780;
wire n10782;
wire n10784;
wire n10785;
wire n10786;
wire n10787;
wire n10788;
wire n10789;
wire n10790;
wire n10792;
wire n10794;
wire n10796;
wire n10798;
wire n10800;
wire n10801;
wire n10803;
wire n10804;
wire n10805;
wire n10807;
wire n10808;
wire n10810;
wire n10811;
wire n10813;
wire n10814;
wire n10815;
wire n10818;
wire n1082;
wire n10820;
wire n10822;
wire n10823;
wire n10824;
wire n10825;
wire n10826;
wire n10827;
wire n10830;
wire n10831;
wire n10833;
wire n10834;
wire n10835;
wire n10836;
wire n10837;
wire n10838;
wire n10839;
wire n10840;
wire n10841;
wire n10842;
wire n10843;
wire n10844;
wire n10845;
wire n10846;
wire n10847;
wire n10848;
wire n10850;
wire n10852;
wire n10853;
wire n10855;
wire n10856;
wire n10857;
wire n10859;
wire n10860;
wire n10861;
wire n10863;
wire n10864;
wire n10865;
wire n10866;
wire n10867;
wire n10868;
wire n1087;
wire n10870;
wire n10871;
wire n10872;
wire n10873;
wire n10874;
wire n10875;
wire n10876;
wire n10877;
wire n10878;
wire n10880;
wire n10881;
wire n10882;
wire n10883;
wire n10884;
wire n10887;
wire n10888;
wire n10890;
wire n10891;
wire n10893;
wire n10894;
wire n10895;
wire n10896;
wire n10897;
wire n10898;
wire n10900;
wire n10902;
wire n10903;
wire n10904;
wire n10905;
wire n10906;
wire n10908;
wire n10909;
wire n10911;
wire n10912;
wire n10913;
wire n10915;
wire n10917;
wire n10918;
wire n10919;
wire n1092;
wire n10920;
wire n10921;
wire n10922;
wire n10924;
wire n10925;
wire n10926;
wire n10927;
wire n10928;
wire n10929;
wire n10932;
wire n10933;
wire n10934;
wire n10936;
wire n10937;
wire n10938;
wire n10940;
wire n10941;
wire n10942;
wire n10943;
wire n10946;
wire n10948;
wire n10949;
wire n10950;
wire n10951;
wire n10952;
wire n10953;
wire n10954;
wire n10955;
wire n10956;
wire n10957;
wire n10958;
wire n10959;
wire n10960;
wire n10961;
wire n10962;
wire n10963;
wire n10964;
wire n10965;
wire n10966;
wire n10967;
wire n10968;
wire n10969;
wire n1097;
wire n10970;
wire n10971;
wire n10972;
wire n10973;
wire n10974;
wire n10975;
wire n10976;
wire n10977;
wire n10978;
wire n10979;
wire n10980;
wire n10981;
wire n10982;
wire n10983;
wire n10984;
wire n10985;
wire n10986;
wire n10987;
wire n10988;
wire n10989;
wire n10990;
wire n10991;
wire n10992;
wire n10993;
wire n10994;
wire n10996;
wire n10997;
wire n10998;
wire n10999;
wire n11000;
wire n11002;
wire n11003;
wire n11004;
wire n11006;
wire n11008;
wire n11009;
wire n11011;
wire n11012;
wire n11013;
wire n11014;
wire n11015;
wire n11016;
wire n11017;
wire n11018;
wire n11019;
wire n1102;
wire n11020;
wire n11024;
wire n11025;
wire n11026;
wire n11029;
wire n11030;
wire n11031;
wire n11033;
wire n11035;
wire n11037;
wire n11038;
wire n11040;
wire n11042;
wire n11043;
wire n11044;
wire n11046;
wire n11047;
wire n11049;
wire n11050;
wire n11052;
wire n11053;
wire n11055;
wire n11056;
wire n11057;
wire n11058;
wire n11059;
wire n11060;
wire n11061;
wire n11062;
wire n11063;
wire n11064;
wire n11065;
wire n11066;
wire n11068;
wire n11069;
wire n1107;
wire n11070;
wire n11072;
wire n11073;
wire n11074;
wire n11077;
wire n11078;
wire n11079;
wire n11081;
wire n11082;
wire n11083;
wire n11084;
wire n11085;
wire n11086;
wire n11088;
wire n11089;
wire n11090;
wire n11091;
wire n11092;
wire n11093;
wire n11094;
wire n11095;
wire n11096;
wire n11098;
wire n11100;
wire n11101;
wire n11102;
wire n11104;
wire n11106;
wire n11107;
wire n11108;
wire n11109;
wire n1111;
wire n11110;
wire n11111;
wire n11112;
wire n11113;
wire n11114;
wire n11115;
wire n11116;
wire n11117;
wire n11118;
wire n11119;
wire n11120;
wire n11121;
wire n11122;
wire n11123;
wire n11125;
wire n11126;
wire n11128;
wire n11130;
wire n11131;
wire n11132;
wire n11133;
wire n11134;
wire n11135;
wire n11136;
wire n11137;
wire n11139;
wire n11140;
wire n11141;
wire n11143;
wire n11145;
wire n11146;
wire n11147;
wire n11148;
wire n11149;
wire n11150;
wire n11151;
wire n11152;
wire n11153;
wire n11155;
wire n11156;
wire n11157;
wire n11158;
wire n11159;
wire n1116;
wire n11160;
wire n11161;
wire n11162;
wire n11163;
wire n11165;
wire n11166;
wire n11167;
wire n11168;
wire n11170;
wire n11172;
wire n11173;
wire n11174;
wire n11175;
wire n11176;
wire n11177;
wire n11178;
wire n11179;
wire n11180;
wire n11182;
wire n11183;
wire n11185;
wire n11186;
wire n11188;
wire n11189;
wire n11191;
wire n11193;
wire n11194;
wire n11196;
wire n11197;
wire n11198;
wire n11200;
wire n11202;
wire n11203;
wire n11204;
wire n11205;
wire n11206;
wire n11207;
wire n11208;
wire n1121;
wire n11210;
wire n11211;
wire n11212;
wire n11213;
wire n11214;
wire n11215;
wire n11216;
wire n11218;
wire n11219;
wire n11220;
wire n11221;
wire n11222;
wire n11223;
wire n11224;
wire n11225;
wire n11226;
wire n11227;
wire n11228;
wire n11229;
wire n11230;
wire n11231;
wire n11232;
wire n11233;
wire n11234;
wire n11235;
wire n11236;
wire n11237;
wire n11238;
wire n11240;
wire n11241;
wire n11243;
wire n11244;
wire n11245;
wire n11246;
wire n11248;
wire n11249;
wire n1125;
wire n11251;
wire n11252;
wire n11254;
wire n11256;
wire n11257;
wire n11258;
wire n11260;
wire n11261;
wire n11262;
wire n11265;
wire n11266;
wire n11267;
wire n11268;
wire n11270;
wire n11271;
wire n11273;
wire n11275;
wire n11276;
wire n11278;
wire n11279;
wire n11281;
wire n11282;
wire n11283;
wire n11286;
wire n11287;
wire n11288;
wire n11289;
wire n11290;
wire n11291;
wire n11292;
wire n11294;
wire n11296;
wire n11297;
wire n11298;
wire n1130;
wire n11300;
wire n11301;
wire n11303;
wire n11305;
wire n11306;
wire n11307;
wire n11308;
wire n11309;
wire n11310;
wire n11311;
wire n11312;
wire n11313;
wire n11314;
wire n11315;
wire n11316;
wire n11317;
wire n11318;
wire n11319;
wire n11320;
wire n11321;
wire n11322;
wire n11323;
wire n11324;
wire n11325;
wire n11326;
wire n11328;
wire n11330;
wire n11331;
wire n11332;
wire n11333;
wire n11334;
wire n11335;
wire n11336;
wire n11337;
wire n11338;
wire n11339;
wire n11340;
wire n11342;
wire n11343;
wire n11345;
wire n11346;
wire n11348;
wire n11349;
wire n1135;
wire n11350;
wire n11352;
wire n11354;
wire n11355;
wire n11356;
wire n11357;
wire n11358;
wire n11359;
wire n11360;
wire n11362;
wire n11363;
wire n11364;
wire n11365;
wire n11366;
wire n11367;
wire n11369;
wire n11370;
wire n11372;
wire n11374;
wire n11375;
wire n11376;
wire n11377;
wire n11378;
wire n11379;
wire n11380;
wire n11381;
wire n11382;
wire n11383;
wire n11384;
wire n11385;
wire n11386;
wire n11387;
wire n11388;
wire n11389;
wire n11390;
wire n11391;
wire n11392;
wire n11393;
wire n11394;
wire n11395;
wire n11396;
wire n11397;
wire n11398;
wire n11399;
wire n1140;
wire n11400;
wire n11401;
wire n11402;
wire n11403;
wire n11404;
wire n11406;
wire n11407;
wire n11408;
wire n11409;
wire n11410;
wire n11411;
wire n11412;
wire n11413;
wire n11414;
wire n11415;
wire n11416;
wire n11417;
wire n11418;
wire n11419;
wire n11420;
wire n11421;
wire n11422;
wire n11423;
wire n11424;
wire n11425;
wire n11426;
wire n11427;
wire n11428;
wire n11429;
wire n11430;
wire n11431;
wire n11432;
wire n11433;
wire n11434;
wire n11435;
wire n11436;
wire n11437;
wire n11439;
wire n11440;
wire n11441;
wire n11442;
wire n11443;
wire n11444;
wire n11445;
wire n11447;
wire n11448;
wire n11449;
wire n1145;
wire n11451;
wire n11452;
wire n11453;
wire n11454;
wire n11455;
wire n11456;
wire n11457;
wire n11458;
wire n11459;
wire n11460;
wire n11461;
wire n11462;
wire n11463;
wire n11464;
wire n11466;
wire n11468;
wire n11469;
wire n11470;
wire n11471;
wire n11472;
wire n11473;
wire n11474;
wire n11475;
wire n11476;
wire n11477;
wire n11478;
wire n11479;
wire n11480;
wire n11481;
wire n11483;
wire n11484;
wire n11485;
wire n11488;
wire n11489;
wire n11490;
wire n11492;
wire n11494;
wire n11495;
wire n11497;
wire n11498;
wire n11499;
wire n1150;
wire n11501;
wire n11502;
wire n11503;
wire n11504;
wire n11506;
wire n11507;
wire n11508;
wire n11509;
wire n11510;
wire n11511;
wire n11512;
wire n11514;
wire n11515;
wire n11516;
wire n11517;
wire n11519;
wire n11520;
wire n11521;
wire n11522;
wire n11523;
wire n11524;
wire n11527;
wire n11528;
wire n11529;
wire n11531;
wire n11533;
wire n11534;
wire n11535;
wire n11536;
wire n11537;
wire n11538;
wire n11539;
wire n11540;
wire n11541;
wire n11542;
wire n11543;
wire n11546;
wire n11547;
wire n11549;
wire n1155;
wire n11551;
wire n11552;
wire n11553;
wire n11554;
wire n11555;
wire n11556;
wire n11557;
wire n11558;
wire n11559;
wire n11560;
wire n11561;
wire n11563;
wire n11564;
wire n11565;
wire n11566;
wire n11567;
wire n11568;
wire n11569;
wire n11571;
wire n11572;
wire n11573;
wire n11574;
wire n11575;
wire n11576;
wire n11577;
wire n11578;
wire n11580;
wire n11581;
wire n11582;
wire n11583;
wire n11584;
wire n11585;
wire n11586;
wire n11587;
wire n11588;
wire n11589;
wire n11590;
wire n11591;
wire n11592;
wire n11593;
wire n11595;
wire n11596;
wire n11597;
wire n11599;
wire n1160;
wire n11600;
wire n11601;
wire n11603;
wire n11604;
wire n11605;
wire n11607;
wire n11608;
wire n11609;
wire n11611;
wire n11612;
wire n11613;
wire n11615;
wire n11616;
wire n11617;
wire n11618;
wire n11619;
wire n11620;
wire n11621;
wire n11622;
wire n11624;
wire n11626;
wire n11627;
wire n11629;
wire n11631;
wire n11633;
wire n11634;
wire n11637;
wire n11638;
wire n11640;
wire n11641;
wire n11642;
wire n11644;
wire n11646;
wire n11647;
wire n11649;
wire n1165;
wire n11650;
wire n11653;
wire n11654;
wire n11655;
wire n11657;
wire n11658;
wire n11659;
wire n11660;
wire n11662;
wire n11663;
wire n11665;
wire n11666;
wire n11667;
wire n11669;
wire n11670;
wire n11672;
wire n11673;
wire n11675;
wire n11676;
wire n11677;
wire n11678;
wire n11679;
wire n11680;
wire n11681;
wire n11682;
wire n11683;
wire n11684;
wire n11685;
wire n11686;
wire n11687;
wire n11688;
wire n11689;
wire n11690;
wire n11692;
wire n11694;
wire n11695;
wire n11696;
wire n11697;
wire n11698;
wire n11699;
wire n1170;
wire n11700;
wire n11701;
wire n11702;
wire n11703;
wire n11704;
wire n11705;
wire n11706;
wire n11707;
wire n11708;
wire n11709;
wire n11710;
wire n11711;
wire n11712;
wire n11713;
wire n11714;
wire n11715;
wire n11716;
wire n11717;
wire n11718;
wire n11719;
wire n11720;
wire n11721;
wire n11722;
wire n11723;
wire n11724;
wire n11725;
wire n11726;
wire n11728;
wire n11729;
wire n11730;
wire n11734;
wire n11735;
wire n11736;
wire n11737;
wire n11738;
wire n11739;
wire n11740;
wire n11741;
wire n11743;
wire n11745;
wire n11746;
wire n11748;
wire n11749;
wire n1175;
wire n11750;
wire n11751;
wire n11752;
wire n11753;
wire n11754;
wire n11755;
wire n11756;
wire n11759;
wire n11760;
wire n11761;
wire n11762;
wire n11763;
wire n11764;
wire n11765;
wire n11767;
wire n11768;
wire n11771;
wire n11773;
wire n11774;
wire n11776;
wire n11777;
wire n11778;
wire n11779;
wire n11780;
wire n11781;
wire n11783;
wire n11786;
wire n11787;
wire n11789;
wire n1179;
wire n11790;
wire n11791;
wire n11793;
wire n11794;
wire n11795;
wire n11796;
wire n11797;
wire n11798;
wire n11799;
wire n11800;
wire n11801;
wire n11803;
wire n11805;
wire n11807;
wire n11808;
wire n11809;
wire n11810;
wire n11811;
wire n11812;
wire n11814;
wire n11815;
wire n11816;
wire n11818;
wire n11820;
wire n11821;
wire n11822;
wire n11823;
wire n11824;
wire n11825;
wire n11828;
wire n11829;
wire n1183;
wire n11830;
wire n11832;
wire n11833;
wire n11835;
wire n11836;
wire n11837;
wire n11838;
wire n11839;
wire n11840;
wire n11841;
wire n11842;
wire n11843;
wire n11844;
wire n11845;
wire n11846;
wire n11847;
wire n11849;
wire n11851;
wire n11852;
wire n11854;
wire n11855;
wire n11856;
wire n11858;
wire n11859;
wire n11860;
wire n11861;
wire n11863;
wire n11864;
wire n11865;
wire n11866;
wire n11868;
wire n11869;
wire n11870;
wire n11872;
wire n11874;
wire n11875;
wire n11877;
wire n11878;
wire n11879;
wire n1188;
wire n11881;
wire n11882;
wire n11884;
wire n11886;
wire n11887;
wire n11888;
wire n11890;
wire n11891;
wire n11893;
wire n11895;
wire n11896;
wire n11898;
wire n11899;
wire n11900;
wire n11902;
wire n11903;
wire n11904;
wire n11905;
wire n11906;
wire n11907;
wire n11909;
wire n11911;
wire n11913;
wire n11914;
wire n11915;
wire n11916;
wire n11917;
wire n11918;
wire n11919;
wire n11920;
wire n11922;
wire n11923;
wire n11924;
wire n11925;
wire n11926;
wire n11927;
wire n11928;
wire n11929;
wire n1193;
wire n11930;
wire n11931;
wire n11932;
wire n11933;
wire n11934;
wire n11935;
wire n11936;
wire n11937;
wire n11938;
wire n11939;
wire n11940;
wire n11941;
wire n11942;
wire n11943;
wire n11944;
wire n11945;
wire n11946;
wire n11947;
wire n11948;
wire n11949;
wire n11950;
wire n11951;
wire n11952;
wire n11953;
wire n11954;
wire n11956;
wire n11957;
wire n11958;
wire n11961;
wire n11962;
wire n11964;
wire n11966;
wire n11968;
wire n11969;
wire n11970;
wire n11971;
wire n11972;
wire n11973;
wire n11974;
wire n11975;
wire n11976;
wire n11977;
wire n11978;
wire n11979;
wire n1198;
wire n11980;
wire n11981;
wire n11982;
wire n11983;
wire n11984;
wire n11985;
wire n11986;
wire n11987;
wire n11988;
wire n11989;
wire n11990;
wire n11991;
wire n11992;
wire n11993;
wire n11995;
wire n11997;
wire n11998;
wire n12000;
wire n12001;
wire n12002;
wire n12004;
wire n12005;
wire n12006;
wire n12008;
wire n12009;
wire n12010;
wire n12011;
wire n12012;
wire n12013;
wire n12014;
wire n12015;
wire n12017;
wire n12018;
wire n12019;
wire n12020;
wire n12021;
wire n12022;
wire n12023;
wire n12025;
wire n12026;
wire n12027;
wire n12029;
wire n1203;
wire n12030;
wire n12032;
wire n12033;
wire n12035;
wire n12036;
wire n12037;
wire n12038;
wire n12039;
wire n12040;
wire n12041;
wire n12042;
wire n12044;
wire n12045;
wire n12046;
wire n12047;
wire n12048;
wire n12049;
wire n12050;
wire n12051;
wire n12053;
wire n12055;
wire n12057;
wire n12058;
wire n12059;
wire n12060;
wire n12061;
wire n12062;
wire n12063;
wire n12064;
wire n12065;
wire n12066;
wire n12067;
wire n12068;
wire n12069;
wire n12070;
wire n12071;
wire n12072;
wire n12073;
wire n12074;
wire n12075;
wire n12076;
wire n12077;
wire n12078;
wire n12079;
wire n1208;
wire n12080;
wire n12081;
wire n12082;
wire n12083;
wire n12084;
wire n12085;
wire n12086;
wire n12087;
wire n12088;
wire n12089;
wire n12091;
wire n12093;
wire n12095;
wire n12096;
wire n12098;
wire n12100;
wire n12101;
wire n12102;
wire n12103;
wire n12104;
wire n12105;
wire n12106;
wire n12108;
wire n12109;
wire n12111;
wire n12112;
wire n12113;
wire n12116;
wire n12118;
wire n12119;
wire n12121;
wire n12122;
wire n12123;
wire n12125;
wire n12127;
wire n12129;
wire n1213;
wire n12130;
wire n12131;
wire n12132;
wire n12134;
wire n12135;
wire n12136;
wire n12138;
wire n12139;
wire n12140;
wire n12142;
wire n12143;
wire n12144;
wire n12145;
wire n12146;
wire n12147;
wire n12148;
wire n12149;
wire n12150;
wire n12151;
wire n12152;
wire n12153;
wire n12154;
wire n12155;
wire n12156;
wire n12158;
wire n12159;
wire n12162;
wire n12163;
wire n12164;
wire n12165;
wire n12166;
wire n12168;
wire n12169;
wire n12170;
wire n12172;
wire n12174;
wire n12175;
wire n12178;
wire n12179;
wire n1218;
wire n12180;
wire n12182;
wire n12183;
wire n12184;
wire n12185;
wire n12186;
wire n12187;
wire n12188;
wire n12189;
wire n12191;
wire n12192;
wire n12193;
wire n12194;
wire n12195;
wire n12196;
wire n12197;
wire n12198;
wire n12199;
wire n12201;
wire n12202;
wire n12204;
wire n12205;
wire n12207;
wire n12208;
wire n12209;
wire n12211;
wire n12212;
wire n12214;
wire n12216;
wire n12217;
wire n12218;
wire n12219;
wire n1222;
wire n12220;
wire n12221;
wire n12222;
wire n12223;
wire n12224;
wire n12225;
wire n12226;
wire n12227;
wire n12228;
wire n12229;
wire n12230;
wire n12231;
wire n12232;
wire n12234;
wire n12235;
wire n12237;
wire n12238;
wire n12239;
wire n12240;
wire n12241;
wire n12242;
wire n12243;
wire n12244;
wire n12245;
wire n12246;
wire n12247;
wire n12248;
wire n12249;
wire n12250;
wire n12251;
wire n12252;
wire n12253;
wire n12254;
wire n12255;
wire n12256;
wire n12257;
wire n12258;
wire n12259;
wire n12260;
wire n12261;
wire n12262;
wire n12263;
wire n12264;
wire n12265;
wire n12266;
wire n12267;
wire n12268;
wire n1227;
wire n12270;
wire n12271;
wire n12273;
wire n12274;
wire n12275;
wire n12276;
wire n12277;
wire n12278;
wire n12279;
wire n12280;
wire n12282;
wire n12283;
wire n12285;
wire n12286;
wire n12287;
wire n12289;
wire n12290;
wire n12291;
wire n12293;
wire n12294;
wire n12295;
wire n12297;
wire n12298;
wire n12299;
wire n12300;
wire n12301;
wire n12302;
wire n12303;
wire n12305;
wire n12307;
wire n12309;
wire n12312;
wire n12313;
wire n12314;
wire n12316;
wire n12318;
wire n12319;
wire n1232;
wire n12320;
wire n12322;
wire n12323;
wire n12324;
wire n12325;
wire n12327;
wire n12329;
wire n12330;
wire n12332;
wire n12333;
wire n12334;
wire n12335;
wire n12336;
wire n12337;
wire n12339;
wire n12341;
wire n12342;
wire n12344;
wire n12345;
wire n12346;
wire n12348;
wire n12349;
wire n12351;
wire n12352;
wire n12354;
wire n12355;
wire n12356;
wire n12358;
wire n12359;
wire n12360;
wire n12361;
wire n12362;
wire n12363;
wire n12364;
wire n12365;
wire n12366;
wire n12367;
wire n12368;
wire n12369;
wire n1237;
wire n12370;
wire n12371;
wire n12372;
wire n12373;
wire n12374;
wire n12375;
wire n12376;
wire n12377;
wire n12378;
wire n12379;
wire n12381;
wire n12382;
wire n12383;
wire n12384;
wire n12385;
wire n12386;
wire n12387;
wire n12388;
wire n12390;
wire n12391;
wire n12392;
wire n12394;
wire n12396;
wire n12397;
wire n12398;
wire n12399;
wire n12401;
wire n12402;
wire n12403;
wire n12404;
wire n12405;
wire n12406;
wire n12407;
wire n12408;
wire n12409;
wire n12410;
wire n12411;
wire n12412;
wire n12413;
wire n12414;
wire n12415;
wire n12416;
wire n12417;
wire n12418;
wire n12419;
wire n1242;
wire n12420;
wire n12421;
wire n12422;
wire n12423;
wire n12424;
wire n12425;
wire n12426;
wire n12427;
wire n12428;
wire n12430;
wire n12431;
wire n12432;
wire n12433;
wire n12434;
wire n12435;
wire n12436;
wire n12437;
wire n12438;
wire n12439;
wire n12440;
wire n12442;
wire n12443;
wire n12444;
wire n12445;
wire n12446;
wire n12448;
wire n12449;
wire n12451;
wire n12452;
wire n12454;
wire n12455;
wire n12456;
wire n12457;
wire n12458;
wire n12459;
wire n12461;
wire n12463;
wire n12464;
wire n12465;
wire n12466;
wire n12467;
wire n12468;
wire n12469;
wire n1247;
wire n12470;
wire n12471;
wire n12472;
wire n12473;
wire n12474;
wire n12475;
wire n12477;
wire n12478;
wire n12480;
wire n12482;
wire n12483;
wire n12486;
wire n12487;
wire n12488;
wire n12490;
wire n12491;
wire n12492;
wire n12493;
wire n12495;
wire n12496;
wire n12498;
wire n12500;
wire n12501;
wire n12502;
wire n12503;
wire n12504;
wire n12505;
wire n12506;
wire n12507;
wire n12508;
wire n12509;
wire n12510;
wire n12511;
wire n12512;
wire n12514;
wire n12515;
wire n12516;
wire n12517;
wire n12518;
wire n12519;
wire n1252;
wire n12520;
wire n12521;
wire n12523;
wire n12525;
wire n12527;
wire n12528;
wire n12529;
wire n12531;
wire n12532;
wire n12533;
wire n12535;
wire n12537;
wire n12538;
wire n12539;
wire n12540;
wire n12541;
wire n12542;
wire n12543;
wire n12545;
wire n12547;
wire n12549;
wire n12550;
wire n12551;
wire n12552;
wire n12553;
wire n12554;
wire n12555;
wire n12556;
wire n12557;
wire n12559;
wire n12560;
wire n12562;
wire n12563;
wire n12565;
wire n12566;
wire n12567;
wire n12569;
wire n1257;
wire n12570;
wire n12571;
wire n12573;
wire n12574;
wire n12576;
wire n12577;
wire n12578;
wire n12579;
wire n12580;
wire n12581;
wire n12583;
wire n12584;
wire n12586;
wire n12587;
wire n12589;
wire n12590;
wire n12592;
wire n12593;
wire n12595;
wire n12598;
wire n12600;
wire n12602;
wire n12603;
wire n12604;
wire n12605;
wire n12606;
wire n12607;
wire n12609;
wire n12610;
wire n12611;
wire n12612;
wire n12613;
wire n12614;
wire n12615;
wire n12616;
wire n12617;
wire n12618;
wire n12619;
wire n1262;
wire n12620;
wire n12621;
wire n12622;
wire n12623;
wire n12624;
wire n12626;
wire n12627;
wire n12628;
wire n12629;
wire n12630;
wire n12632;
wire n12634;
wire n12635;
wire n12636;
wire n12638;
wire n12639;
wire n12640;
wire n12641;
wire n12642;
wire n12643;
wire n12644;
wire n12645;
wire n12646;
wire n12647;
wire n12648;
wire n12650;
wire n12651;
wire n12652;
wire n12653;
wire n12654;
wire n12655;
wire n12656;
wire n12657;
wire n12658;
wire n12660;
wire n12661;
wire n12662;
wire n12663;
wire n12664;
wire n12666;
wire n12668;
wire n12669;
wire n1267;
wire n12671;
wire n12672;
wire n12673;
wire n12676;
wire n12677;
wire n12679;
wire n12681;
wire n12682;
wire n12683;
wire n12685;
wire n12686;
wire n12687;
wire n12688;
wire n12689;
wire n12690;
wire n12691;
wire n12692;
wire n12693;
wire n12695;
wire n12696;
wire n12697;
wire n12700;
wire n12701;
wire n12702;
wire n12703;
wire n12704;
wire n12705;
wire n12706;
wire n12707;
wire n12708;
wire n12710;
wire n12711;
wire n12712;
wire n12714;
wire n12715;
wire n12716;
wire n12717;
wire n12719;
wire n1272;
wire n12720;
wire n12721;
wire n12722;
wire n12723;
wire n12724;
wire n12726;
wire n12727;
wire n12728;
wire n12729;
wire n12730;
wire n12731;
wire n12732;
wire n12733;
wire n12734;
wire n12735;
wire n12736;
wire n12737;
wire n12738;
wire n12739;
wire n12741;
wire n12742;
wire n12743;
wire n12746;
wire n12748;
wire n12749;
wire n12750;
wire n12751;
wire n12752;
wire n12753;
wire n12755;
wire n12756;
wire n12757;
wire n12759;
wire n12761;
wire n12762;
wire n12763;
wire n12765;
wire n12767;
wire n12768;
wire n1277;
wire n12770;
wire n12771;
wire n12773;
wire n12774;
wire n12775;
wire n12777;
wire n12778;
wire n12780;
wire n12781;
wire n12782;
wire n12783;
wire n12785;
wire n12786;
wire n12788;
wire n12789;
wire n12790;
wire n12791;
wire n12792;
wire n12793;
wire n12794;
wire n12797;
wire n12798;
wire n12799;
wire n12801;
wire n12802;
wire n12803;
wire n12804;
wire n12805;
wire n12806;
wire n12807;
wire n12808;
wire n12809;
wire n12810;
wire n12811;
wire n12814;
wire n12815;
wire n12817;
wire n12819;
wire n1282;
wire n12820;
wire n12821;
wire n12822;
wire n12823;
wire n12824;
wire n12826;
wire n12827;
wire n12829;
wire n12830;
wire n12831;
wire n12832;
wire n12835;
wire n12836;
wire n12837;
wire n12838;
wire n12839;
wire n12840;
wire n12841;
wire n12842;
wire n12843;
wire n12844;
wire n12845;
wire n12846;
wire n12847;
wire n12848;
wire n12849;
wire n12850;
wire n12851;
wire n12852;
wire n12853;
wire n12854;
wire n12855;
wire n12856;
wire n12857;
wire n12858;
wire n12859;
wire n1286;
wire n12860;
wire n12862;
wire n12863;
wire n12865;
wire n12866;
wire n12867;
wire n12869;
wire n12870;
wire n12872;
wire n12873;
wire n12874;
wire n12875;
wire n12876;
wire n12878;
wire n12879;
wire n12880;
wire n12881;
wire n12883;
wire n12884;
wire n12885;
wire n12886;
wire n12888;
wire n12889;
wire n12890;
wire n12892;
wire n12894;
wire n12895;
wire n12896;
wire n12897;
wire n12898;
wire n12899;
wire n12900;
wire n12901;
wire n12903;
wire n12904;
wire n12905;
wire n12906;
wire n12907;
wire n12908;
wire n1291;
wire n12910;
wire n12911;
wire n12913;
wire n12914;
wire n12915;
wire n12918;
wire n12919;
wire n12920;
wire n12922;
wire n12923;
wire n12925;
wire n12926;
wire n12927;
wire n12929;
wire n12930;
wire n12931;
wire n12933;
wire n12934;
wire n12935;
wire n12936;
wire n12937;
wire n12938;
wire n12939;
wire n12940;
wire n12941;
wire n12942;
wire n12943;
wire n12945;
wire n12946;
wire n12948;
wire n12949;
wire n12951;
wire n12953;
wire n12954;
wire n12955;
wire n12957;
wire n12958;
wire n12959;
wire n1296;
wire n12960;
wire n12961;
wire n12963;
wire n12965;
wire n12966;
wire n12967;
wire n12968;
wire n12969;
wire n12970;
wire n12971;
wire n12972;
wire n12973;
wire n12975;
wire n12976;
wire n12977;
wire n12978;
wire n12979;
wire n12980;
wire n12981;
wire n12982;
wire n12984;
wire n12985;
wire n12986;
wire n12988;
wire n12989;
wire n12990;
wire n12993;
wire n12996;
wire n12997;
wire n12999;
wire n13002;
wire n13003;
wire n13004;
wire n13006;
wire n13007;
wire n1301;
wire n13011;
wire n13012;
wire n13013;
wire n13014;
wire n13015;
wire n13016;
wire n13017;
wire n13019;
wire n13020;
wire n13021;
wire n13022;
wire n13023;
wire n13024;
wire n13025;
wire n13026;
wire n13028;
wire n13029;
wire n13030;
wire n13032;
wire n13033;
wire n13035;
wire n13036;
wire n13039;
wire n13040;
wire n13043;
wire n13044;
wire n13046;
wire n13047;
wire n13049;
wire n13050;
wire n13051;
wire n13052;
wire n13053;
wire n13054;
wire n13055;
wire n13056;
wire n13057;
wire n13058;
wire n1306;
wire n13060;
wire n13061;
wire n13062;
wire n13063;
wire n13064;
wire n13065;
wire n13066;
wire n13067;
wire n13068;
wire n13069;
wire n13070;
wire n13071;
wire n13072;
wire n13073;
wire n13074;
wire n13076;
wire n13077;
wire n13079;
wire n13080;
wire n13082;
wire n13083;
wire n13085;
wire n13086;
wire n13087;
wire n13089;
wire n13092;
wire n13093;
wire n13094;
wire n13096;
wire n13097;
wire n13098;
wire n13099;
wire n1310;
wire n13101;
wire n13102;
wire n13104;
wire n13105;
wire n13106;
wire n13107;
wire n13108;
wire n13109;
wire n13110;
wire n13111;
wire n13112;
wire n13113;
wire n13114;
wire n13115;
wire n13116;
wire n13119;
wire n13120;
wire n13121;
wire n13122;
wire n13123;
wire n13126;
wire n13127;
wire n13128;
wire n13129;
wire n13130;
wire n13131;
wire n13132;
wire n13133;
wire n13134;
wire n13136;
wire n13137;
wire n13138;
wire n13139;
wire n13140;
wire n13142;
wire n13143;
wire n13144;
wire n13145;
wire n13146;
wire n13147;
wire n13148;
wire n13149;
wire n1315;
wire n13150;
wire n13151;
wire n13152;
wire n13153;
wire n13154;
wire n13155;
wire n13157;
wire n13158;
wire n13160;
wire n13161;
wire n13162;
wire n13164;
wire n13165;
wire n13167;
wire n13168;
wire n13170;
wire n13172;
wire n13173;
wire n13175;
wire n13176;
wire n13179;
wire n13180;
wire n13182;
wire n13183;
wire n13185;
wire n13186;
wire n13187;
wire n13189;
wire n13191;
wire n13193;
wire n13195;
wire n13196;
wire n13198;
wire n1320;
wire n13200;
wire n13201;
wire n13203;
wire n13204;
wire n13206;
wire n13207;
wire n13209;
wire n13210;
wire n13211;
wire n13212;
wire n13213;
wire n13214;
wire n13215;
wire n13216;
wire n13217;
wire n13218;
wire n13219;
wire n13220;
wire n13222;
wire n13224;
wire n13225;
wire n13226;
wire n13227;
wire n13228;
wire n13229;
wire n13230;
wire n13232;
wire n13234;
wire n13236;
wire n13237;
wire n13238;
wire n13240;
wire n13241;
wire n13242;
wire n13243;
wire n13244;
wire n13245;
wire n13246;
wire n13247;
wire n13248;
wire n13249;
wire n1325;
wire n13250;
wire n13251;
wire n13253;
wire n13254;
wire n13255;
wire n13257;
wire n13258;
wire n13259;
wire n13261;
wire n13263;
wire n13264;
wire n13265;
wire n13267;
wire n13268;
wire n13270;
wire n13271;
wire n13272;
wire n13273;
wire n13274;
wire n13275;
wire n13276;
wire n13277;
wire n13278;
wire n13279;
wire n13280;
wire n13281;
wire n13282;
wire n13283;
wire n13284;
wire n13286;
wire n13287;
wire n13288;
wire n13290;
wire n13291;
wire n13292;
wire n13293;
wire n13294;
wire n13295;
wire n13296;
wire n13297;
wire n13298;
wire n13299;
wire n1330;
wire n13300;
wire n13301;
wire n13303;
wire n13304;
wire n13306;
wire n13307;
wire n13308;
wire n13310;
wire n13311;
wire n13312;
wire n13314;
wire n13316;
wire n13317;
wire n13318;
wire n13320;
wire n13322;
wire n13324;
wire n13325;
wire n13326;
wire n13327;
wire n13328;
wire n13329;
wire n13330;
wire n13331;
wire n13332;
wire n13333;
wire n13335;
wire n13336;
wire n13337;
wire n13339;
wire n13340;
wire n13341;
wire n13342;
wire n13343;
wire n13344;
wire n13345;
wire n13346;
wire n13347;
wire n13348;
wire n13349;
wire n1335;
wire n13350;
wire n13351;
wire n13352;
wire n13353;
wire n13354;
wire n13356;
wire n13358;
wire n13359;
wire n13360;
wire n13361;
wire n13364;
wire n13365;
wire n13366;
wire n13368;
wire n13369;
wire n13371;
wire n13372;
wire n13373;
wire n13374;
wire n13375;
wire n13376;
wire n13377;
wire n13378;
wire n13380;
wire n13381;
wire n13383;
wire n13384;
wire n13385;
wire n13386;
wire n13387;
wire n13388;
wire n13389;
wire n1339;
wire n13390;
wire n13391;
wire n13392;
wire n13393;
wire n13395;
wire n13396;
wire n13397;
wire n13398;
wire n13399;
wire n13400;
wire n13401;
wire n13402;
wire n13403;
wire n13405;
wire n13406;
wire n13409;
wire n13411;
wire n13412;
wire n13413;
wire n13414;
wire n13415;
wire n13416;
wire n13417;
wire n13418;
wire n13419;
wire n13420;
wire n13421;
wire n13422;
wire n13424;
wire n13426;
wire n13427;
wire n13428;
wire n13429;
wire n13430;
wire n13431;
wire n13432;
wire n13434;
wire n13435;
wire n13436;
wire n13437;
wire n13438;
wire n13439;
wire n1344;
wire n13440;
wire n13441;
wire n13442;
wire n13443;
wire n13444;
wire n13445;
wire n13446;
wire n13447;
wire n13448;
wire n13449;
wire n13450;
wire n13451;
wire n13452;
wire n13453;
wire n13454;
wire n13455;
wire n13456;
wire n13457;
wire n13458;
wire n13459;
wire n13460;
wire n13461;
wire n13462;
wire n13463;
wire n13464;
wire n13465;
wire n13467;
wire n13468;
wire n13470;
wire n13471;
wire n13472;
wire n13473;
wire n13475;
wire n13476;
wire n13477;
wire n13480;
wire n13482;
wire n13484;
wire n13485;
wire n13486;
wire n13488;
wire n1349;
wire n13490;
wire n13491;
wire n13492;
wire n13493;
wire n13494;
wire n13495;
wire n13496;
wire n13497;
wire n13498;
wire n13499;
wire n13500;
wire n13501;
wire n13502;
wire n13503;
wire n13504;
wire n13505;
wire n13506;
wire n13507;
wire n13508;
wire n13509;
wire n13510;
wire n13511;
wire n13512;
wire n13513;
wire n13514;
wire n13515;
wire n13516;
wire n13517;
wire n13518;
wire n13519;
wire n13520;
wire n13521;
wire n13522;
wire n13523;
wire n13524;
wire n13525;
wire n13526;
wire n13527;
wire n13529;
wire n13530;
wire n13531;
wire n13533;
wire n13535;
wire n13536;
wire n13537;
wire n13539;
wire n1354;
wire n13540;
wire n13542;
wire n13543;
wire n13544;
wire n13546;
wire n13547;
wire n13548;
wire n13550;
wire n13551;
wire n13552;
wire n13554;
wire n13555;
wire n13556;
wire n13558;
wire n13559;
wire n13560;
wire n13562;
wire n13566;
wire n13567;
wire n13569;
wire n13571;
wire n13572;
wire n13573;
wire n13575;
wire n13576;
wire n13577;
wire n13578;
wire n13579;
wire n13581;
wire n13582;
wire n13583;
wire n13585;
wire n13586;
wire n13589;
wire n1359;
wire n13590;
wire n13591;
wire n13592;
wire n13593;
wire n13594;
wire n13595;
wire n13596;
wire n13598;
wire n13600;
wire n13601;
wire n13602;
wire n13603;
wire n13604;
wire n13605;
wire n13606;
wire n13607;
wire n13609;
wire n13610;
wire n13612;
wire n13613;
wire n13616;
wire n13619;
wire n13620;
wire n13621;
wire n13623;
wire n13624;
wire n13625;
wire n13627;
wire n13629;
wire n13630;
wire n13631;
wire n13632;
wire n13634;
wire n13635;
wire n13637;
wire n13638;
wire n13639;
wire n1364;
wire n13640;
wire n13641;
wire n13642;
wire n13643;
wire n13645;
wire n13646;
wire n13647;
wire n13648;
wire n13649;
wire n13650;
wire n13651;
wire n13652;
wire n13654;
wire n13655;
wire n13656;
wire n13657;
wire n13658;
wire n13659;
wire n13660;
wire n13661;
wire n13662;
wire n13663;
wire n13664;
wire n13665;
wire n13666;
wire n13668;
wire n13670;
wire n13671;
wire n13673;
wire n13674;
wire n13675;
wire n13676;
wire n13677;
wire n13678;
wire n13679;
wire n13680;
wire n13682;
wire n13683;
wire n13685;
wire n13687;
wire n13689;
wire n1369;
wire n13690;
wire n13691;
wire n13693;
wire n13695;
wire n13697;
wire n13699;
wire n13701;
wire n13702;
wire n13704;
wire n13706;
wire n13708;
wire n13709;
wire n13711;
wire n13712;
wire n13714;
wire n13715;
wire n13719;
wire n13721;
wire n13722;
wire n13723;
wire n13726;
wire n13727;
wire n13728;
wire n13730;
wire n13732;
wire n13734;
wire n13735;
wire n13737;
wire n13738;
wire n13739;
wire n1374;
wire n13740;
wire n13742;
wire n13743;
wire n13745;
wire n13746;
wire n13748;
wire n13749;
wire n13751;
wire n13752;
wire n13753;
wire n13754;
wire n13755;
wire n13756;
wire n13757;
wire n13758;
wire n13760;
wire n13761;
wire n13762;
wire n13763;
wire n13764;
wire n13765;
wire n13767;
wire n13768;
wire n13769;
wire n13770;
wire n13771;
wire n13772;
wire n13773;
wire n13774;
wire n13775;
wire n13776;
wire n13777;
wire n13778;
wire n13779;
wire n13780;
wire n13782;
wire n13784;
wire n13787;
wire n13788;
wire n1379;
wire n13790;
wire n13792;
wire n13793;
wire n13795;
wire n13797;
wire n13799;
wire n13801;
wire n13802;
wire n13804;
wire n13805;
wire n13806;
wire n13807;
wire n13808;
wire n13809;
wire n13810;
wire n13811;
wire n13812;
wire n13813;
wire n13814;
wire n13815;
wire n13816;
wire n13817;
wire n13818;
wire n13819;
wire n13820;
wire n13822;
wire n13824;
wire n13825;
wire n13826;
wire n13828;
wire n13829;
wire n13830;
wire n13833;
wire n13835;
wire n13836;
wire n13837;
wire n13839;
wire n1384;
wire n13841;
wire n13842;
wire n13843;
wire n13845;
wire n13846;
wire n13847;
wire n13849;
wire n13850;
wire n13851;
wire n13853;
wire n13854;
wire n13856;
wire n13857;
wire n13858;
wire n13860;
wire n13862;
wire n13863;
wire n13864;
wire n13865;
wire n13867;
wire n13869;
wire n13871;
wire n13872;
wire n13873;
wire n13875;
wire n13877;
wire n13878;
wire n13879;
wire n1388;
wire n13881;
wire n13883;
wire n13884;
wire n13885;
wire n13886;
wire n13887;
wire n13888;
wire n13890;
wire n13891;
wire n13892;
wire n13895;
wire n13896;
wire n13897;
wire n13901;
wire n13902;
wire n13903;
wire n13905;
wire n13906;
wire n13908;
wire n13909;
wire n13910;
wire n13912;
wire n13913;
wire n13914;
wire n13916;
wire n13917;
wire n13919;
wire n1392;
wire n13920;
wire n13922;
wire n13923;
wire n13924;
wire n13926;
wire n13927;
wire n13928;
wire n13929;
wire n13930;
wire n13931;
wire n13932;
wire n13933;
wire n13934;
wire n13935;
wire n13937;
wire n13938;
wire n13940;
wire n13941;
wire n13942;
wire n13944;
wire n13946;
wire n13947;
wire n13948;
wire n13950;
wire n13951;
wire n13953;
wire n13954;
wire n13955;
wire n13956;
wire n13957;
wire n13958;
wire n13959;
wire n13961;
wire n13964;
wire n13965;
wire n13966;
wire n13968;
wire n13969;
wire n1397;
wire n13970;
wire n13971;
wire n13973;
wire n13975;
wire n13976;
wire n13978;
wire n13979;
wire n13981;
wire n13982;
wire n13984;
wire n13986;
wire n13988;
wire n13989;
wire n13990;
wire n13991;
wire n13992;
wire n13993;
wire n13994;
wire n13995;
wire n13996;
wire n13997;
wire n13998;
wire n13999;
wire n14000;
wire n14001;
wire n14002;
wire n14003;
wire n14004;
wire n14006;
wire n14007;
wire n14008;
wire n14009;
wire n1401;
wire n14010;
wire n14011;
wire n14013;
wire n14014;
wire n14015;
wire n14016;
wire n14017;
wire n14018;
wire n14019;
wire n14021;
wire n14022;
wire n14024;
wire n14025;
wire n14026;
wire n14027;
wire n14028;
wire n14029;
wire n14030;
wire n14031;
wire n14033;
wire n14034;
wire n14035;
wire n14036;
wire n14037;
wire n14038;
wire n14039;
wire n14040;
wire n14041;
wire n14042;
wire n14043;
wire n14045;
wire n14046;
wire n14048;
wire n14049;
wire n14050;
wire n14052;
wire n14053;
wire n14054;
wire n14057;
wire n14058;
wire n14059;
wire n1406;
wire n14061;
wire n14062;
wire n14064;
wire n14066;
wire n14068;
wire n14069;
wire n14071;
wire n14072;
wire n14074;
wire n14075;
wire n14077;
wire n14078;
wire n14079;
wire n14080;
wire n14081;
wire n14082;
wire n14083;
wire n14084;
wire n14087;
wire n14088;
wire n14091;
wire n14092;
wire n14094;
wire n14096;
wire n14097;
wire n14100;
wire n14101;
wire n14102;
wire n14104;
wire n14105;
wire n14106;
wire n14107;
wire n14108;
wire n14109;
wire n1411;
wire n14111;
wire n14113;
wire n14114;
wire n14115;
wire n14116;
wire n14117;
wire n14118;
wire n14119;
wire n14120;
wire n14121;
wire n14123;
wire n14125;
wire n14127;
wire n14128;
wire n14130;
wire n14131;
wire n14132;
wire n14133;
wire n14134;
wire n14137;
wire n14139;
wire n14140;
wire n14141;
wire n14142;
wire n14143;
wire n14144;
wire n14145;
wire n14146;
wire n14147;
wire n14148;
wire n14149;
wire n1415;
wire n14150;
wire n14151;
wire n14153;
wire n14154;
wire n14157;
wire n14158;
wire n14160;
wire n14161;
wire n14162;
wire n14163;
wire n14165;
wire n14166;
wire n14167;
wire n14168;
wire n14169;
wire n14170;
wire n14171;
wire n14173;
wire n14175;
wire n14176;
wire n14177;
wire n14178;
wire n14179;
wire n14180;
wire n14181;
wire n14182;
wire n14183;
wire n14184;
wire n14185;
wire n14186;
wire n14187;
wire n14188;
wire n14189;
wire n14190;
wire n14191;
wire n14193;
wire n14195;
wire n14196;
wire n14198;
wire n14199;
wire n1420;
wire n14201;
wire n14202;
wire n14203;
wire n14204;
wire n14205;
wire n14208;
wire n14209;
wire n14211;
wire n14212;
wire n14213;
wire n14215;
wire n14216;
wire n14218;
wire n14219;
wire n14220;
wire n14221;
wire n14222;
wire n14223;
wire n14224;
wire n14225;
wire n14226;
wire n14227;
wire n14228;
wire n14229;
wire n14230;
wire n14231;
wire n14232;
wire n14234;
wire n14235;
wire n14238;
wire n14239;
wire n14240;
wire n14241;
wire n14242;
wire n14243;
wire n14244;
wire n14245;
wire n14246;
wire n14247;
wire n14248;
wire n14249;
wire n1425;
wire n14250;
wire n14252;
wire n14254;
wire n14255;
wire n14256;
wire n14259;
wire n14260;
wire n14261;
wire n14262;
wire n14263;
wire n14264;
wire n14266;
wire n14267;
wire n14269;
wire n14270;
wire n14271;
wire n14273;
wire n14274;
wire n14275;
wire n14276;
wire n14277;
wire n14279;
wire n14281;
wire n14282;
wire n14283;
wire n14285;
wire n14286;
wire n14287;
wire n14288;
wire n14289;
wire n14290;
wire n14291;
wire n14292;
wire n14293;
wire n14294;
wire n14295;
wire n14296;
wire n14297;
wire n14298;
wire n14299;
wire n1430;
wire n14300;
wire n14301;
wire n14302;
wire n14303;
wire n14304;
wire n14305;
wire n14306;
wire n14309;
wire n14310;
wire n14314;
wire n14315;
wire n14316;
wire n14317;
wire n14318;
wire n14319;
wire n14320;
wire n14321;
wire n14322;
wire n14323;
wire n14324;
wire n14326;
wire n14327;
wire n14328;
wire n14329;
wire n14330;
wire n14331;
wire n14333;
wire n14334;
wire n14336;
wire n14337;
wire n14338;
wire n14339;
wire n14340;
wire n14341;
wire n14343;
wire n14344;
wire n14345;
wire n14346;
wire n14347;
wire n14348;
wire n14349;
wire n1435;
wire n14350;
wire n14352;
wire n14353;
wire n14355;
wire n14356;
wire n14357;
wire n14359;
wire n14360;
wire n14361;
wire n14363;
wire n14364;
wire n14365;
wire n14366;
wire n14367;
wire n14368;
wire n14370;
wire n14371;
wire n14372;
wire n14376;
wire n14377;
wire n14378;
wire n14379;
wire n14380;
wire n14381;
wire n14382;
wire n14383;
wire n14384;
wire n14385;
wire n14386;
wire n14387;
wire n14388;
wire n14389;
wire n14391;
wire n14392;
wire n14394;
wire n14398;
wire n14399;
wire n1440;
wire n14401;
wire n14403;
wire n14404;
wire n14405;
wire n14406;
wire n14408;
wire n14409;
wire n14411;
wire n14412;
wire n14414;
wire n14415;
wire n14417;
wire n14419;
wire n14420;
wire n14422;
wire n14423;
wire n14425;
wire n14426;
wire n14427;
wire n14429;
wire n14431;
wire n14432;
wire n14433;
wire n14435;
wire n14436;
wire n14438;
wire n14439;
wire n1444;
wire n14441;
wire n14442;
wire n14443;
wire n14444;
wire n14446;
wire n14447;
wire n14448;
wire n14449;
wire n14450;
wire n14451;
wire n14452;
wire n14454;
wire n14455;
wire n14456;
wire n14457;
wire n14458;
wire n14459;
wire n14460;
wire n14461;
wire n14462;
wire n14463;
wire n14464;
wire n14465;
wire n14466;
wire n14467;
wire n14468;
wire n14469;
wire n14470;
wire n14471;
wire n14472;
wire n14473;
wire n14474;
wire n14475;
wire n14476;
wire n14477;
wire n14478;
wire n14479;
wire n14480;
wire n14481;
wire n14482;
wire n14483;
wire n14484;
wire n14485;
wire n14486;
wire n14488;
wire n14489;
wire n1449;
wire n14490;
wire n14491;
wire n14492;
wire n14493;
wire n14494;
wire n14495;
wire n14496;
wire n14497;
wire n14498;
wire n14499;
wire n14500;
wire n14502;
wire n14503;
wire n14504;
wire n14505;
wire n14506;
wire n14507;
wire n14508;
wire n14509;
wire n14510;
wire n14511;
wire n14513;
wire n14514;
wire n14516;
wire n14518;
wire n14519;
wire n14521;
wire n14523;
wire n14524;
wire n14526;
wire n14527;
wire n14529;
wire n14530;
wire n14531;
wire n14533;
wire n14535;
wire n14538;
wire n14539;
wire n1454;
wire n14540;
wire n14541;
wire n14542;
wire n14543;
wire n14544;
wire n14545;
wire n14547;
wire n14548;
wire n14549;
wire n14551;
wire n14552;
wire n14556;
wire n14558;
wire n14559;
wire n14560;
wire n14561;
wire n14563;
wire n14564;
wire n14565;
wire n14566;
wire n14567;
wire n14569;
wire n14571;
wire n14572;
wire n14574;
wire n14575;
wire n14577;
wire n14578;
wire n14580;
wire n14581;
wire n14585;
wire n14586;
wire n14588;
wire n14589;
wire n1459;
wire n14590;
wire n14592;
wire n14593;
wire n14594;
wire n14597;
wire n14599;
wire n14602;
wire n14603;
wire n14604;
wire n14606;
wire n14607;
wire n14609;
wire n14611;
wire n14612;
wire n14614;
wire n14615;
wire n14616;
wire n14617;
wire n14620;
wire n14621;
wire n14622;
wire n14623;
wire n14625;
wire n14626;
wire n14627;
wire n14628;
wire n14629;
wire n14630;
wire n14631;
wire n14632;
wire n14633;
wire n14634;
wire n14635;
wire n14636;
wire n14637;
wire n14638;
wire n14639;
wire n1464;
wire n14640;
wire n14641;
wire n14642;
wire n14643;
wire n14644;
wire n14645;
wire n14646;
wire n14647;
wire n14648;
wire n14649;
wire n14650;
wire n14651;
wire n14652;
wire n14653;
wire n14654;
wire n14655;
wire n14656;
wire n14658;
wire n14659;
wire n14660;
wire n14661;
wire n14662;
wire n14664;
wire n14665;
wire n14666;
wire n14669;
wire n14670;
wire n14672;
wire n14673;
wire n14674;
wire n14677;
wire n14679;
wire n14680;
wire n14681;
wire n14682;
wire n14683;
wire n14684;
wire n14685;
wire n14687;
wire n14688;
wire n14689;
wire n1469;
wire n14690;
wire n14691;
wire n14693;
wire n14695;
wire n14696;
wire n14697;
wire n14698;
wire n14699;
wire n14700;
wire n14701;
wire n14702;
wire n14703;
wire n14704;
wire n14705;
wire n14706;
wire n14708;
wire n14709;
wire n14710;
wire n14712;
wire n14713;
wire n14714;
wire n14715;
wire n14717;
wire n14718;
wire n14719;
wire n14720;
wire n14721;
wire n14723;
wire n14724;
wire n14725;
wire n14726;
wire n14727;
wire n14729;
wire n14730;
wire n14731;
wire n14732;
wire n14733;
wire n14734;
wire n14736;
wire n14737;
wire n14739;
wire n1474;
wire n14740;
wire n14741;
wire n14742;
wire n14743;
wire n14744;
wire n14745;
wire n14746;
wire n14748;
wire n14750;
wire n14751;
wire n14752;
wire n14754;
wire n14756;
wire n14757;
wire n14759;
wire n14760;
wire n14761;
wire n14762;
wire n14763;
wire n14764;
wire n14765;
wire n14766;
wire n14767;
wire n14768;
wire n14769;
wire n14771;
wire n14772;
wire n14775;
wire n14776;
wire n14778;
wire n14779;
wire n1478;
wire n14780;
wire n14782;
wire n14783;
wire n14784;
wire n14786;
wire n14787;
wire n14789;
wire n14791;
wire n14792;
wire n14793;
wire n14795;
wire n14798;
wire n14799;
wire n14801;
wire n14803;
wire n14804;
wire n14806;
wire n14807;
wire n14808;
wire n14810;
wire n14812;
wire n14814;
wire n14816;
wire n14817;
wire n14819;
wire n14820;
wire n14821;
wire n14822;
wire n14823;
wire n14824;
wire n14826;
wire n14828;
wire n14829;
wire n1483;
wire n14830;
wire n14831;
wire n14832;
wire n14833;
wire n14834;
wire n14836;
wire n14837;
wire n14838;
wire n14840;
wire n14841;
wire n14842;
wire n14843;
wire n14844;
wire n14845;
wire n14846;
wire n14847;
wire n14848;
wire n14849;
wire n14850;
wire n14851;
wire n14852;
wire n14853;
wire n14854;
wire n14855;
wire n14856;
wire n14857;
wire n14859;
wire n14860;
wire n14861;
wire n14862;
wire n14864;
wire n14865;
wire n14866;
wire n14867;
wire n14868;
wire n14869;
wire n14870;
wire n14871;
wire n14872;
wire n14873;
wire n14874;
wire n14875;
wire n14876;
wire n14877;
wire n14878;
wire n14879;
wire n1488;
wire n14880;
wire n14881;
wire n14882;
wire n14883;
wire n14884;
wire n14885;
wire n14886;
wire n14887;
wire n14888;
wire n14889;
wire n14890;
wire n14891;
wire n14892;
wire n14893;
wire n14894;
wire n14895;
wire n14896;
wire n14898;
wire n14899;
wire n14902;
wire n14903;
wire n14904;
wire n14905;
wire n14906;
wire n14907;
wire n14908;
wire n14909;
wire n14910;
wire n14911;
wire n14912;
wire n14913;
wire n14914;
wire n14915;
wire n14916;
wire n14918;
wire n14919;
wire n1492;
wire n14920;
wire n14921;
wire n14922;
wire n14923;
wire n14924;
wire n14925;
wire n14926;
wire n14928;
wire n14929;
wire n14930;
wire n14931;
wire n14932;
wire n14933;
wire n14934;
wire n14935;
wire n14937;
wire n14938;
wire n14939;
wire n14940;
wire n14941;
wire n14942;
wire n14943;
wire n14944;
wire n14946;
wire n14947;
wire n14948;
wire n14950;
wire n14951;
wire n14953;
wire n14955;
wire n14956;
wire n14958;
wire n14959;
wire n14962;
wire n14963;
wire n14964;
wire n14965;
wire n14966;
wire n14967;
wire n14968;
wire n14969;
wire n1497;
wire n14970;
wire n14972;
wire n14973;
wire n14974;
wire n14975;
wire n14976;
wire n14977;
wire n14979;
wire n14980;
wire n14982;
wire n14984;
wire n14985;
wire n14986;
wire n14987;
wire n14988;
wire n14989;
wire n14990;
wire n14991;
wire n14992;
wire n14994;
wire n14996;
wire n14997;
wire n14998;
wire n15000;
wire n15001;
wire n15002;
wire n15003;
wire n15004;
wire n15005;
wire n15006;
wire n15007;
wire n15008;
wire n15010;
wire n15011;
wire n15012;
wire n15013;
wire n15014;
wire n15015;
wire n15016;
wire n15017;
wire n15018;
wire n15019;
wire n1502;
wire n15020;
wire n15021;
wire n15022;
wire n15023;
wire n15024;
wire n15025;
wire n15026;
wire n15028;
wire n15029;
wire n15030;
wire n15032;
wire n15034;
wire n15035;
wire n15036;
wire n15037;
wire n15039;
wire n15040;
wire n15041;
wire n15043;
wire n15044;
wire n15046;
wire n15047;
wire n15048;
wire n15049;
wire n15054;
wire n15055;
wire n15056;
wire n15057;
wire n15058;
wire n15060;
wire n15061;
wire n15063;
wire n15065;
wire n15066;
wire n15067;
wire n15068;
wire n15069;
wire n1507;
wire n15070;
wire n15071;
wire n15072;
wire n15074;
wire n1512;
wire n1517;
wire n1521;
wire n1526;
wire n1531;
wire n1536;
wire n1540;
wire n1545;
wire n1549;
wire n1554;
wire n1559;
wire n1564;
wire n1569;
wire n1574;
wire n1579;
wire n1582;
wire n1587;
wire n1592;
wire n1597;
wire n1602;
wire n1605;
wire n1609;
wire n1614;
wire n1618;
wire n1623;
wire n1627;
wire n1631;
wire n1636;
wire n1641;
wire n1646;
wire n1651;
wire n1656;
wire n1661;
wire n1666;
wire n1671;
wire n1676;
wire n1681;
wire n1686;
wire n1691;
wire n1696;
wire n1701;
wire n1706;
wire n1711;
wire n1715;
wire n1720;
wire n1725;
wire n1730;
wire n1735;
wire n1739;
wire n1744;
wire n1749;
wire n1754;
wire n1759;
wire n1764;
wire n1769;
wire n1774;
wire n1779;
wire n1783;
wire n1787;
wire n1792;
wire n1797;
wire n1802;
wire n1807;
wire n1812;
wire n1817;
wire n1822;
wire n1826;
wire n1831;
wire n1835;
wire n1839;
wire n1844;
wire n1849;
wire n1854;
wire n1859;
wire n1863;
wire n1868;
wire n1872;
wire n1877;
wire n1881;
wire n1886;
wire n1891;
wire n1896;
wire n1901;
wire n1906;
wire n1911;
wire n1916;
wire n1921;
wire n1926;
wire n1931;
wire n1936;
wire n1941;
wire n1946;
wire n1951;
wire n1956;
wire n1960;
wire n1965;
wire n1970;
wire n1975;
wire n1980;
wire n1985;
wire n1990;
wire n1995;
wire n2000;
wire n2005;
wire n2010;
wire n2015;
wire n2020;
wire n2025;
wire n2030;
wire n2035;
wire n2040;
wire n2045;
wire n2050;
wire n2055;
wire n2060;
wire n2065;
wire n2070;
wire n2075;
wire n2080;
wire n2085;
wire n2090;
wire n2095;
wire n2100;
wire n2105;
wire n2110;
wire n2115;
wire n2120;
wire n2125;
wire n2130;
wire n2135;
wire n2140;
wire n2145;
wire n2150;
wire n2155;
wire n2160;
wire n2165;
wire n2169;
wire n2174;
wire n2179;
wire n2184;
wire n2189;
wire n2193;
wire n2198;
wire n2202;
wire n2207;
wire n2212;
wire n2217;
wire n2222;
wire n2227;
wire n2232;
wire n2237;
wire n2242;
wire n2246;
wire n2251;
wire n2256;
wire n2261;
wire n2266;
wire n2271;
wire n2276;
wire n2281;
wire n2286;
wire n2291;
wire n2296;
wire n2301;
wire n2306;
wire n2311;
wire n2316;
wire n2321;
wire n2325;
wire n2330;
wire n2334;
wire n2338;
wire n2342;
wire n2347;
wire n2352;
wire n2357;
wire n2362;
wire n2367;
wire n2371;
wire n2375;
wire n2380;
wire n2385;
wire n2390;
wire n2395;
wire n2400;
wire n2404;
wire n2409;
wire n2414;
wire n2419;
wire n2424;
wire n2429;
wire n2434;
wire n2439;
wire n2444;
wire n2449;
wire n2453;
wire n2458;
wire n2463;
wire n2468;
wire n2473;
wire n2477;
wire n2482;
wire n2487;
wire n2492;
wire n2497;
wire n2502;
wire n2507;
wire n2512;
wire n2517;
wire n2522;
wire n2527;
wire n2532;
wire n2537;
wire n2541;
wire n2546;
wire n2551;
wire n2556;
wire n2560;
wire n2564;
wire n2568;
wire n2572;
wire n2577;
wire n2582;
wire n2587;
wire n2592;
wire n2597;
wire n2602;
wire n2607;
wire n2612;
wire n2617;
wire n2622;
wire n2627;
wire n2632;
wire n2637;
wire n2642;
wire n2647;
wire n2652;
wire n2657;
wire n2662;
wire n2667;
wire n2671;
wire n2676;
wire n2681;
wire n2685;
wire n2690;
wire n2695;
wire n2700;
wire n2705;
wire n2710;
wire n2715;
wire n2720;
wire n2725;
wire n2730;
wire n2735;
wire n2740;
wire n2745;
wire n2750;
wire n2755;
wire n2760;
wire n2765;
wire n2769;
wire n2774;
wire n2779;
wire n2784;
wire n2789;
wire n2794;
wire n2798;
wire n2803;
wire n2808;
wire n2813;
wire n2817;
wire n2822;
wire n2827;
wire n2832;
wire n2836;
wire n2841;
wire n2846;
wire n2851;
wire n2855;
wire n2860;
wire n2864;
wire n2869;
wire n2874;
wire n2878;
wire n2883;
wire n2888;
wire n2893;
wire n2898;
wire n2903;
wire n2908;
wire n2912;
wire n2917;
wire n2922;
wire n2927;
wire n2932;
wire n2937;
wire n2942;
wire n2946;
wire n2951;
wire n2956;
wire n2960;
wire n2965;
wire n2970;
wire n2975;
wire n2980;
wire n2985;
wire n2990;
wire n2995;
wire n3000;
wire n3005;
wire n3010;
wire n3015;
wire n3020;
wire n3025;
wire n3030;
wire n3034;
wire n3039;
wire n3043;
wire n3048;
wire n3053;
wire n3058;
wire n3063;
wire n3068;
wire n3073;
wire n3077;
wire n3082;
wire n3087;
wire n3092;
wire n3097;
wire n3101;
wire n3106;
wire n3111;
wire n3116;
wire n3121;
wire n3126;
wire n3131;
wire n3136;
wire n3141;
wire n3146;
wire n3151;
wire n3156;
wire n3161;
wire n3166;
wire n3171;
wire n3176;
wire n3181;
wire n3186;
wire n3191;
wire n3195;
wire n3200;
wire n3205;
wire n3210;
wire n3215;
wire n3220;
wire n3225;
wire n3230;
wire n3234;
wire n3238;
wire n3243;
wire n3247;
wire n3252;
wire n3257;
wire n3262;
wire n3267;
wire n3272;
wire n3277;
wire n3282;
wire n3287;
wire n3291;
wire n3296;
wire n3300;
wire n3305;
wire n3310;
wire n3315;
wire n3320;
wire n3325;
wire n3330;
wire n3335;
wire n3340;
wire n3345;
wire n3350;
wire n3355;
wire n3359;
wire n3364;
wire n3369;
wire n3374;
wire n3379;
wire n3384;
wire n3389;
wire n3394;
wire n3399;
wire n3404;
wire n3409;
wire n3413;
wire n3416;
wire n3421;
wire n3426;
wire n3430;
wire n3435;
wire n3440;
wire n3445;
wire n3450;
wire n3455;
wire n3460;
wire n3465;
wire n3470;
wire n3475;
wire n3480;
wire n3485;
wire n3490;
wire n3495;
wire n3499;
wire n3504;
wire n3509;
wire n3513;
wire n3518;
wire n3523;
wire n3528;
wire n3533;
wire n3538;
wire n3543;
wire n3548;
wire n3553;
wire n3558;
wire n3563;
wire n3568;
wire n3573;
wire n3578;
wire n3583;
wire n3588;
wire n3593;
wire n3598;
wire n3603;
wire n3608;
wire n3613;
wire n3618;
wire n3623;
wire n3628;
wire n3633;
wire n3638;
wire n3642;
wire n3647;
wire n3652;
wire n3657;
wire n3662;
wire n3667;
wire n3672;
wire n3677;
wire n3682;
wire n3687;
wire n3692;
wire n3697;
wire n3702;
wire n3707;
wire n3712;
wire n3717;
wire n3722;
wire n3727;
wire n3732;
wire n3737;
wire n3742;
wire n3746;
wire n3750;
wire n3754;
wire n3758;
wire n3763;
wire n3768;
wire n3773;
wire n3778;
wire n3782;
wire n3787;
wire n3792;
wire n3796;
wire n3801;
wire n3805;
wire n3810;
wire n3815;
wire n3820;
wire n3825;
wire n3830;
wire n3835;
wire n3839;
wire n3844;
wire n3849;
wire n3854;
wire n3859;
wire n3864;
wire n3869;
wire n3874;
wire n3879;
wire n3884;
wire n3889;
wire n3894;
wire n3899;
wire n3904;
wire n3909;
wire n3914;
wire n3919;
wire n3923;
wire n3928;
wire n3933;
wire n3937;
wire n3942;
wire n3947;
wire n3952;
wire n3957;
wire n3962;
wire n3967;
wire n3972;
wire n3976;
wire n3980;
wire n3985;
wire n3990;
wire n3994;
wire n3999;
wire n4004;
wire n4009;
wire n4014;
wire n4019;
wire n4024;
wire n4029;
wire n4034;
wire n4039;
wire n4044;
wire n4049;
wire n4054;
wire n4059;
wire n4064;
wire n4069;
wire n4074;
wire n4079;
wire n4084;
wire n4088;
wire n4093;
wire n4098;
wire n4103;
wire n4108;
wire n4112;
wire n4116;
wire n4120;
wire n4124;
wire n4129;
wire n4133;
wire n4137;
wire n4142;
wire n4147;
wire n4151;
wire n4156;
wire n4161;
wire n4165;
wire n4170;
wire n4175;
wire n4180;
wire n4185;
wire n4190;
wire n4195;
wire n4200;
wire n4205;
wire n4210;
wire n4215;
wire n4220;
wire n4225;
wire n4230;
wire n4235;
wire n4240;
wire n4245;
wire n4250;
wire n4255;
wire n4259;
wire n4264;
wire n4269;
wire n4274;
wire n4279;
wire n4283;
wire n4288;
wire n4293;
wire n4298;
wire n4303;
wire n4308;
wire n4312;
wire n4316;
wire n4321;
wire n4326;
wire n4331;
wire n4336;
wire n4341;
wire n4346;
wire n4351;
wire n4355;
wire n4360;
wire n4364;
wire n4368;
wire n4372;
wire n4377;
wire n4382;
wire n4387;
wire n4392;
wire n4397;
wire n4401;
wire n4405;
wire n4410;
wire n4415;
wire n4420;
wire n4425;
wire n4430;
wire n4434;
wire n4439;
wire n4444;
wire n4449;
wire n4454;
wire n4459;
wire n4463;
wire n4468;
wire n4473;
wire n4477;
wire n4482;
wire n4487;
wire n4491;
wire n4496;
wire n4501;
wire n4506;
wire n4511;
wire n4516;
wire n4521;
wire n4525;
wire n4530;
wire n4535;
wire n4539;
wire n4544;
wire n4549;
wire n4554;
wire n4559;
wire n4564;
wire n4569;
wire n4574;
wire n4579;
wire n4584;
wire n4589;
wire n4594;
wire n4598;
wire n4603;
wire n4608;
wire n4613;
wire n4618;
wire n4623;
wire n4627;
wire n4632;
wire n4637;
wire n4642;
wire n4647;
wire n4650;
wire n4654;
wire n4659;
wire n4664;
wire n4668;
wire n4673;
wire n4678;
wire n4682;
wire n4687;
wire n4692;
wire n4696;
wire n4700;
wire n4705;
wire n4710;
wire n4715;
wire n4719;
wire n4724;
wire n4729;
wire n4734;
wire n4739;
wire n4744;
wire n4749;
wire n4754;
wire n4759;
wire n4764;
wire n4769;
wire n4774;
wire n4779;
wire n4784;
wire n4788;
wire n4793;
wire n4797;
wire n4802;
wire n4807;
wire n4812;
wire n4817;
wire n4822;
wire n4827;
wire n4832;
wire n4837;
wire n4842;
wire n4846;
wire n4851;
wire n4856;
wire n4861;
wire n4866;
wire n4871;
wire n4875;
wire n4879;
wire n4884;
wire n4889;
wire n4894;
wire n4899;
wire n4904;
wire n4908;
wire n4913;
wire n4918;
wire n4923;
wire n4927;
wire n4932;
wire n4937;
wire n4941;
wire n4946;
wire n4951;
wire n4956;
wire n4961;
wire n4966;
wire n4971;
wire n4976;
wire n4980;
wire n4985;
wire n4990;
wire n4995;
wire n500;
wire n5000;
wire n5005;
wire n5010;
wire n5015;
wire n5020;
wire n5025;
wire n5030;
wire n5035;
wire n5038;
wire n5043;
wire n5048;
wire n505;
wire n5052;
wire n5057;
wire n5062;
wire n5067;
wire n5072;
wire n5077;
wire n5082;
wire n5087;
wire n5091;
wire n5096;
wire n510;
wire n5101;
wire n5105;
wire n5110;
wire n5115;
wire n5120;
wire n5125;
wire n5130;
wire n5135;
wire n5139;
wire n514;
wire n5143;
wire n5147;
wire n5152;
wire n5157;
wire n5161;
wire n5165;
wire n5169;
wire n5174;
wire n5179;
wire n5184;
wire n5189;
wire n519;
wire n5194;
wire n5198;
wire n5203;
wire n5208;
wire n5212;
wire n5217;
wire n5222;
wire n5227;
wire n5232;
wire n5237;
wire n524;
wire n5242;
wire n5247;
wire n5252;
wire n5257;
wire n5262;
wire n5266;
wire n5270;
wire n5275;
wire n5279;
wire n528;
wire n5283;
wire n5288;
wire n5293;
wire n5297;
wire n5302;
wire n5306;
wire n5311;
wire n5316;
wire n5321;
wire n5326;
wire n533;
wire n5331;
wire n5336;
wire n5341;
wire n5346;
wire n5351;
wire n5355;
wire n5360;
wire n5365;
wire n5370;
wire n5375;
wire n5379;
wire n538;
wire n5384;
wire n5389;
wire n5394;
wire n5399;
wire n5403;
wire n5408;
wire n5412;
wire n5417;
wire n5422;
wire n5427;
wire n543;
wire n5431;
wire n5436;
wire n5441;
wire n5445;
wire n5449;
wire n5454;
wire n5459;
wire n5464;
wire n5469;
wire n5473;
wire n5477;
wire n548;
wire n5481;
wire n5486;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5495_1;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5500_1;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5504_1;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5513;
wire n5513_1;
wire n5514;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5522;
wire n5523;
wire n5523_1;
wire n5525;
wire n5526;
wire n5528;
wire n5528_1;
wire n5529;
wire n553;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5537;
wire n5537_1;
wire n5538;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5546;
wire n5547;
wire n5547_1;
wire n5549;
wire n5550;
wire n5552;
wire n5552_1;
wire n5553;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5561;
wire n5562;
wire n5562_1;
wire n5564;
wire n5565;
wire n5567;
wire n5567_1;
wire n5568;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5576;
wire n5577;
wire n5577_1;
wire n5579;
wire n558;
wire n5580;
wire n5582;
wire n5582_1;
wire n5583;
wire n5585;
wire n5585_1;
wire n5586;
wire n5588;
wire n5589;
wire n5589_1;
wire n5591;
wire n5592;
wire n5594;
wire n5594_1;
wire n5595;
wire n5597;
wire n5597_1;
wire n5598;
wire n5600;
wire n5601;
wire n5601_1;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5609;
wire n5610;
wire n5610_1;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5618;
wire n5619;
wire n5619_1;
wire n5621;
wire n5622;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5629_1;
wire n563;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5637;
wire n5638;
wire n5638_1;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5646;
wire n5647;
wire n5647_1;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5655;
wire n5656;
wire n5656_1;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5661_1;
wire n5662;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5666_1;
wire n5667;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5671_1;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5676_1;
wire n5677;
wire n5678;
wire n5679;
wire n568;
wire n5680;
wire n5681;
wire n5681_1;
wire n5682;
wire n5684;
wire n5685;
wire n5685_1;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5690_1;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5700_1;
wire n5701;
wire n5702;
wire n5703;
wire n5705;
wire n5705_1;
wire n5706;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5710_1;
wire n5711;
wire n5712;
wire n5713;
wire n5714;
wire n5714_1;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5719_1;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5724_1;
wire n5725;
wire n5726;
wire n5727;
wire n5728;
wire n5729;
wire n5729_1;
wire n573;
wire n5730;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5734_1;
wire n5735;
wire n5737;
wire n5738;
wire n5739;
wire n5739_1;
wire n5740;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5744_1;
wire n5746;
wire n5747;
wire n5748;
wire n5748_1;
wire n5749;
wire n5750;
wire n5751;
wire n5752;
wire n5753;
wire n5753_1;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5758_1;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5763_1;
wire n5764;
wire n5766;
wire n5767;
wire n5768;
wire n5768_1;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5773_1;
wire n5774;
wire n5775;
wire n5777;
wire n5777_1;
wire n5778;
wire n5779;
wire n578;
wire n5780;
wire n5781;
wire n5782;
wire n5782_1;
wire n5783;
wire n5784;
wire n5785;
wire n5786;
wire n5787;
wire n5787_1;
wire n5788;
wire n5789;
wire n5790;
wire n5791;
wire n5792;
wire n5792_1;
wire n5793;
wire n5794;
wire n5796;
wire n5797;
wire n5797_1;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5802_1;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5807_1;
wire n5808;
wire n5809;
wire n5811;
wire n5812;
wire n5812_1;
wire n5813;
wire n5814;
wire n5815;
wire n5815_1;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5820_1;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5825;
wire n5826;
wire n5827;
wire n5828;
wire n5829;
wire n583;
wire n5830;
wire n5830_1;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5835;
wire n5835_1;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5839_1;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5844_1;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5849_1;
wire n5850;
wire n5851;
wire n5853;
wire n5853_1;
wire n5854;
wire n5855;
wire n5856;
wire n5857;
wire n5858;
wire n5858_1;
wire n5859;
wire n5860;
wire n5861;
wire n5862;
wire n5863;
wire n5863_1;
wire n5864;
wire n5865;
wire n5866;
wire n5867;
wire n5868;
wire n5868_1;
wire n5869;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5873_1;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5878_1;
wire n5879;
wire n588;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5883_1;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5888_1;
wire n5889;
wire n5890;
wire n5891;
wire n5892;
wire n5893;
wire n5893_1;
wire n5895;
wire n5897;
wire n5898;
wire n5898_1;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5903_1;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5914;
wire n5916;
wire n5917;
wire n5917_1;
wire n5918;
wire n5919;
wire n5920;
wire n5921;
wire n5921_1;
wire n5922;
wire n5923;
wire n5924;
wire n5925;
wire n5926;
wire n5926_1;
wire n5927;
wire n5928;
wire n5929;
wire n593;
wire n5930;
wire n5931;
wire n5931_1;
wire n5932;
wire n5933;
wire n5934;
wire n5935;
wire n5935_1;
wire n5936;
wire n5937;
wire n5938;
wire n5939;
wire n5939_1;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5944;
wire n5944_1;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5949;
wire n5949_1;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5954;
wire n5954_1;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5959;
wire n5959_1;
wire n5960;
wire n5961;
wire n5962;
wire n5963;
wire n5964;
wire n5964_1;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5969;
wire n5969_1;
wire n5970;
wire n5971;
wire n5972;
wire n5973;
wire n5974;
wire n5974_1;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5978_1;
wire n5979;
wire n598;
wire n5980;
wire n5981;
wire n5982;
wire n5983;
wire n5983_1;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5988;
wire n5988_1;
wire n5989;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5993_1;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n5998_1;
wire n5999;
wire n6000;
wire n6001;
wire n6001_1;
wire n6002;
wire n6003;
wire n6004;
wire n6005;
wire n6005_1;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6009_1;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6013_1;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6018_1;
wire n6019;
wire n6020;
wire n6021;
wire n6022;
wire n6023;
wire n6023_1;
wire n6024;
wire n6025;
wire n6026;
wire n6027;
wire n6028;
wire n6028_1;
wire n6029;
wire n603;
wire n6031;
wire n6032;
wire n6033;
wire n6033_1;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6037_1;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6042_1;
wire n6043;
wire n6044;
wire n6045;
wire n6047;
wire n6047_1;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6052_1;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6057_1;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6062_1;
wire n6063;
wire n6065;
wire n6066;
wire n6067;
wire n6067_1;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6072_1;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6077_1;
wire n6078;
wire n6079;
wire n608;
wire n6080;
wire n6081;
wire n6082;
wire n6082_1;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6087_1;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6091_1;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6095_1;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6099_1;
wire n6100;
wire n6101;
wire n6102;
wire n6102_1;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6107_1;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6111_1;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6116_1;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6121_1;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6126_1;
wire n6127;
wire n6128;
wire n6129;
wire n613;
wire n6130;
wire n6131;
wire n6131_1;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6136_1;
wire n6137;
wire n6139;
wire n6140;
wire n6141;
wire n6141_1;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6145_1;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6150_1;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6155_1;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6160_1;
wire n6161;
wire n6163;
wire n6164;
wire n6164_1;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6169_1;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6173_1;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6177_1;
wire n6178;
wire n6179;
wire n618;
wire n6180;
wire n6181;
wire n6181_1;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6186_1;
wire n6187;
wire n6188;
wire n6190;
wire n6191;
wire n6191_1;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6196_1;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6201_1;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6206_1;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6211_1;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6216_1;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6221_1;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6226_1;
wire n6227;
wire n6228;
wire n6229;
wire n623;
wire n6230;
wire n6231;
wire n6231_1;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6235_1;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6240_1;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6244_1;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6249_1;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6254_1;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6258_1;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6263_1;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6268_1;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6272_1;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6277_1;
wire n6278;
wire n6279;
wire n628;
wire n6280;
wire n6281;
wire n6282;
wire n6282_1;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6287_1;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6292_1;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6297_1;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6302_1;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6306_1;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6311_1;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6316_1;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6321_1;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6326_1;
wire n6327;
wire n6328;
wire n6329;
wire n633;
wire n6330;
wire n6331;
wire n6331_1;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6336_1;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6341_1;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6346_1;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6351_1;
wire n6352;
wire n6354;
wire n6355;
wire n6356;
wire n6356_1;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6360_1;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6364_1;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6369_1;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6373_1;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6378_1;
wire n6379;
wire n638;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6383_1;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6388_1;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6393_1;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6397_1;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6401_1;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6406_1;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6411_1;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6416_1;
wire n6417;
wire n6418;
wire n6419;
wire n642;
wire n6420;
wire n6421;
wire n6421_1;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6426_1;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6431_1;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6436_1;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6441_1;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6446_1;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6451_1;
wire n6452;
wire n6454;
wire n6455;
wire n6456;
wire n6456_1;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6460_1;
wire n6461;
wire n6463;
wire n6464;
wire n6464_1;
wire n6465;
wire n6467;
wire n6468;
wire n6469;
wire n6469_1;
wire n647;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6474_1;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6479_1;
wire n6480;
wire n6481;
wire n6483;
wire n6484;
wire n6484_1;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6489_1;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6493_1;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6498_1;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6503_1;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6507_1;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6512_1;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6517_1;
wire n6518;
wire n6519;
wire n652;
wire n6520;
wire n6521;
wire n6522;
wire n6522_1;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6526_1;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6531_1;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6536_1;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6541_1;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6546_1;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6551_1;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6556_1;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6561_1;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6566_1;
wire n6567;
wire n6568;
wire n6569;
wire n657;
wire n6570;
wire n6571;
wire n6571_1;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6575_1;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n6579_1;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6584_1;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6589_1;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6594_1;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6599_1;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6604_1;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6609_1;
wire n661;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6614_1;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6619_1;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6624_1;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6629_1;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6634_1;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6639_1;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6644_1;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6649_1;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6654_1;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6659_1;
wire n666;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6664_1;
wire n6665;
wire n6667;
wire n6668;
wire n6669;
wire n6669_1;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6674_1;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6679_1;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6684_1;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6689_1;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6694_1;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6699_1;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6704_1;
wire n6705;
wire n6707;
wire n6708;
wire n6709;
wire n671;
wire n6711;
wire n6713;
wire n6713_1;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6718_1;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6723_1;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6728_1;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6733_1;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6738_1;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6743_1;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6748_1;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6753_1;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6758_1;
wire n6759;
wire n676;
wire n6760;
wire n6761;
wire n6763;
wire n6763_1;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6773_1;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6778_1;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6782_1;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6786_1;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6791_1;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6796_1;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6801_1;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6806_1;
wire n6807;
wire n6808;
wire n6809;
wire n681;
wire n6810;
wire n6811;
wire n6811_1;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6816_1;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6821_1;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6826_1;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6831;
wire n6831_1;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6836_1;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6841_1;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6846_1;
wire n6847;
wire n6848;
wire n6850;
wire n6851;
wire n6851_1;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6856;
wire n6856_1;
wire n6857;
wire n6858;
wire n6859;
wire n686;
wire n6860;
wire n6861;
wire n6861_1;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6865_1;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6875_1;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n6880;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6885_1;
wire n6886;
wire n6887;
wire n6888;
wire n6890;
wire n6890_1;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6899;
wire n6900;
wire n6900_1;
wire n6902;
wire n6903;
wire n6904;
wire n6905;
wire n6905_1;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n691;
wire n6910;
wire n6910_1;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6914_1;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6919_1;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6924_1;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6929_1;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6934_1;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6939_1;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6944_1;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6949_1;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6954_1;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6958_1;
wire n6959;
wire n696;
wire n6960;
wire n6961;
wire n6962;
wire n6962_1;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6966_1;
wire n6967;
wire n6968;
wire n6970;
wire n6971;
wire n6971_1;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6976_1;
wire n6977;
wire n6979;
wire n6980;
wire n6981;
wire n6981_1;
wire n6983;
wire n6985;
wire n6985_1;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6989_1;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6998_1;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7003_1;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7007_1;
wire n7008;
wire n7009;
wire n701;
wire n7010;
wire n7011;
wire n7012;
wire n7012_1;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7017_1;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7021_1;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7026_1;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7030_1;
wire n7031;
wire n7032;
wire n7033;
wire n7034;
wire n7034_1;
wire n7035;
wire n7036;
wire n7037;
wire n7038;
wire n7039;
wire n7039_1;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7044_1;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7048_1;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7053_1;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7058_1;
wire n7059;
wire n706;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7063_1;
wire n7064;
wire n7065;
wire n7066;
wire n7067;
wire n7068;
wire n7068_1;
wire n7069;
wire n7071;
wire n7072;
wire n7073;
wire n7073_1;
wire n7074;
wire n7075;
wire n7077;
wire n7078;
wire n7078_1;
wire n7080;
wire n7081;
wire n7082;
wire n7082_1;
wire n7084;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7091_1;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7095_1;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7100_1;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7104_1;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7108_1;
wire n7109;
wire n711;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7113_1;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7118_1;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7123_1;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7128_1;
wire n7129;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7133_1;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7138_1;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7143_1;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7148_1;
wire n7149;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7153_1;
wire n7154;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7158_1;
wire n7159;
wire n716;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7163_1;
wire n7164;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7168_1;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7173_1;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7177_1;
wire n7178;
wire n7179;
wire n7180;
wire n7181;
wire n7182;
wire n7182_1;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7187_1;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7192_1;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7197_1;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7202_1;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7206_1;
wire n7207;
wire n7208;
wire n7209;
wire n721;
wire n7210;
wire n7211;
wire n7211_1;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7216_1;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7221_1;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7226_1;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7231_1;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7235_1;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7240_1;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7245;
wire n7245_1;
wire n7246;
wire n7247;
wire n7248;
wire n7249;
wire n7250;
wire n7250_1;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7255_1;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n726;
wire n7260;
wire n7260_1;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7265_1;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n7270;
wire n7270_1;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7275_1;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7280_1;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7285_1;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7290_1;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7295_1;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7300_1;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7304_1;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7308_1;
wire n7309;
wire n731;
wire n7310;
wire n7311;
wire n7312;
wire n7312_1;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7317_1;
wire n7318;
wire n7319;
wire n7320;
wire n7321;
wire n7321_1;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7326_1;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7331_1;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7336_1;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7341;
wire n7341_1;
wire n7342;
wire n7343;
wire n7345;
wire n7346;
wire n7346_1;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7351_1;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7355_1;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n736;
wire n7360;
wire n7361;
wire n7362;
wire n7364;
wire n7365;
wire n7365_1;
wire n7366;
wire n7367;
wire n7369;
wire n7370;
wire n7370_1;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7375_1;
wire n7376;
wire n7377;
wire n7378;
wire n7379;
wire n7379_1;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7384_1;
wire n7385;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7389_1;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7394_1;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7398_1;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7403_1;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7408_1;
wire n7409;
wire n741;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7413_1;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7418_1;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7423_1;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7428_1;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7432_1;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7436_1;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7441_1;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7446_1;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7451_1;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7459;
wire n746;
wire n7460;
wire n7460_1;
wire n7461;
wire n7463;
wire n7464;
wire n7465;
wire n7465_1;
wire n7466;
wire n7467;
wire n7469;
wire n7470;
wire n7470_1;
wire n7471;
wire n7473;
wire n7474;
wire n7475;
wire n7475_1;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7480_1;
wire n7482;
wire n7483;
wire n7484;
wire n7484_1;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7489_1;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7494_1;
wire n7495;
wire n7496;
wire n7497;
wire n7499;
wire n7499_1;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7504_1;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7509_1;
wire n751;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7514_1;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7519_1;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7524_1;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7529_1;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7534_1;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7538_1;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7543_1;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7548_1;
wire n7549;
wire n755;
wire n7550;
wire n7551;
wire n7552;
wire n7552_1;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7557_1;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7562_1;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7566_1;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7571_1;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7575_1;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7580_1;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7585_1;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7590_1;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7595_1;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n760;
wire n7600;
wire n7600_1;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7605_1;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7609_1;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7613_1;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7617_1;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7621_1;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7626_1;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7631_1;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7636_1;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7640_1;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7645_1;
wire n7647;
wire n7648;
wire n765;
wire n7650;
wire n7650_1;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7655;
wire n7655_1;
wire n7657;
wire n7658;
wire n7660;
wire n7660_1;
wire n7661;
wire n7663;
wire n7664;
wire n7665;
wire n7665_1;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7670_1;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7675_1;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7685_1;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7694;
wire n7695;
wire n7695_1;
wire n7696;
wire n7698;
wire n7699;
wire n770;
wire n7700;
wire n7700_1;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7704_1;
wire n7705;
wire n7706;
wire n7708;
wire n7709;
wire n7709_1;
wire n7712;
wire n7713;
wire n7714;
wire n7714_1;
wire n7716;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7724_1;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7734_1;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7738_1;
wire n774;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7743_1;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7748_1;
wire n7750;
wire n7751;
wire n7753;
wire n7753_1;
wire n7754;
wire n7755;
wire n7756;
wire n7758;
wire n7758_1;
wire n7759;
wire n7761;
wire n7762;
wire n7763;
wire n7763_1;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7768_1;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7773_1;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7778_1;
wire n7779;
wire n778;
wire n7780;
wire n7781;
wire n7782;
wire n7782_1;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7787_1;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7792_1;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7796_1;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7801_1;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7806_1;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7811_1;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7816_1;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7821_1;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7826_1;
wire n7827;
wire n7829;
wire n783;
wire n7830;
wire n7830_1;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7834_1;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7843_1;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7848_1;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7853_1;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7857_1;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7862_1;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7870;
wire n7871;
wire n7871_1;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7876_1;
wire n7877;
wire n7878;
wire n7879;
wire n788;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7885_1;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7889_1;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7893_1;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7898_1;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7902_1;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7906_1;
wire n7907;
wire n7908;
wire n7910;
wire n7911;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7916_1;
wire n7917;
wire n7919;
wire n7920;
wire n7921;
wire n7921_1;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7925_1;
wire n7926;
wire n7928;
wire n7929;
wire n793;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7935_1;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7940_1;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7950;
wire n7950_1;
wire n7951;
wire n7952;
wire n7954;
wire n7954_1;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7962_1;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7967_1;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7972_1;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7977_1;
wire n7978;
wire n7979;
wire n798;
wire n7980;
wire n7981;
wire n7982;
wire n7982_1;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7987_1;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7992_1;
wire n7994;
wire n7995;
wire n7996;
wire n7996_1;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8001_1;
wire n8002;
wire n8003;
wire n8004;
wire n8006;
wire n8006_1;
wire n8007;
wire n8008;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8021_1;
wire n8022;
wire n8024;
wire n8025;
wire n8026;
wire n8026_1;
wire n8027;
wire n8028;
wire n8029;
wire n803;
wire n8030;
wire n8031;
wire n8031_1;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8038;
wire n8039;
wire n8041;
wire n8041_1;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8046_1;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8051_1;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8055_1;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8059_1;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8063_1;
wire n8065;
wire n8066;
wire n8067;
wire n8067_1;
wire n8068;
wire n8069;
wire n8071;
wire n8072;
wire n8072_1;
wire n8074;
wire n8075;
wire n8076;
wire n8076_1;
wire n8077;
wire n8078;
wire n8079;
wire n808;
wire n8080;
wire n8081;
wire n8081_1;
wire n8082;
wire n8083;
wire n8085;
wire n8086;
wire n8086_1;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
wire n8091_1;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8101;
wire n8101_1;
wire n8102;
wire n8104;
wire n8105;
wire n8106;
wire n8106_1;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8111_1;
wire n8112;
wire n8114;
wire n8115;
wire n8116;
wire n8116_1;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8125;
wire n8125_1;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n813;
wire n8130;
wire n8130_1;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8135_1;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8140_1;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8145_1;
wire n8146;
wire n8147;
wire n8148;
wire n8150;
wire n8150_1;
wire n8151;
wire n8153;
wire n8155;
wire n8155_1;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8160_1;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8165_1;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8170_1;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8175_1;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n818;
wire n8180;
wire n8180_1;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8185_1;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8190_1;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8195_1;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8200_1;
wire n8201;
wire n8202;
wire n8203;
wire n8205;
wire n8205_1;
wire n8206;
wire n8207;
wire n8209;
wire n8210;
wire n8210_1;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8214_1;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8219_1;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8223_1;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8227_1;
wire n8228;
wire n8229;
wire n823;
wire n8230;
wire n8231;
wire n8231_1;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8235_1;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8240_1;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8245_1;
wire n8246;
wire n8248;
wire n8250;
wire n8250_1;
wire n8251;
wire n8252;
wire n8254;
wire n8255;
wire n8255_1;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8260_1;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8264_1;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8268_1;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8272_1;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8276_1;
wire n8277;
wire n8278;
wire n8279;
wire n828;
wire n8280;
wire n8281;
wire n8282;
wire n8284;
wire n8285;
wire n8286;
wire n8286_1;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8291_1;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8296_1;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8301_1;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8305_1;
wire n8307;
wire n8308;
wire n8310;
wire n8310_1;
wire n8312;
wire n8313;
wire n8315;
wire n8315_1;
wire n8316;
wire n8317;
wire n8319;
wire n8320;
wire n8320_1;
wire n8321;
wire n8322;
wire n8324;
wire n8325;
wire n8325_1;
wire n8326;
wire n8327;
wire n8329;
wire n833;
wire n8330;
wire n8330_1;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8335_1;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8339_1;
wire n8340;
wire n8341;
wire n8342;
wire n8344;
wire n8344_1;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8349_1;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8363;
wire n8363_1;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8372_1;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8376_1;
wire n8377;
wire n8378;
wire n8379;
wire n838;
wire n8380;
wire n8380_1;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8389;
wire n8389_1;
wire n8391;
wire n8392;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8398;
wire n8399;
wire n8399_1;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8404_1;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8409_1;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8414_1;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8424_1;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n8429_1;
wire n843;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8433_1;
wire n8435;
wire n8436;
wire n8437;
wire n8438;
wire n8438_1;
wire n8440;
wire n8442;
wire n8443;
wire n8443_1;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8452_1;
wire n8453;
wire n8454;
wire n8456;
wire n8457;
wire n8457_1;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8462_1;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8467_1;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8472_1;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8477_1;
wire n8478;
wire n8479;
wire n848;
wire n8480;
wire n8481;
wire n8482;
wire n8482_1;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8486_1;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8491_1;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8501_1;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8505_1;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8510_1;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8523;
wire n8524;
wire n8524_1;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8529_1;
wire n853;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8534;
wire n8534_1;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8538_1;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8543_1;
wire n8544;
wire n8546;
wire n8547;
wire n8548;
wire n8548_1;
wire n8550;
wire n8551;
wire n8553;
wire n8553_1;
wire n8554;
wire n8555;
wire n8557;
wire n8558;
wire n8558_1;
wire n8560;
wire n8562;
wire n8562_1;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8567_1;
wire n8568;
wire n8569;
wire n8570;
wire n8572;
wire n8572_1;
wire n8573;
wire n8575;
wire n8576;
wire n8577;
wire n8577_1;
wire n8578;
wire n8579;
wire n858;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8587_1;
wire n8588;
wire n8590;
wire n8592;
wire n8592_1;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8597_1;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8602_1;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8607_1;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8612_1;
wire n8613;
wire n8616;
wire n8616_1;
wire n8617;
wire n8618;
wire n8620;
wire n8621;
wire n8621_1;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n863;
wire n8630;
wire n8631;
wire n8631_1;
wire n8633;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8641_1;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8646_1;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8650_1;
wire n8651;
wire n8652;
wire n8653;
wire n8655;
wire n8655_1;
wire n8656;
wire n8658;
wire n8659;
wire n8659_1;
wire n8661;
wire n8663;
wire n8664;
wire n8664_1;
wire n8665;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8671;
wire n8673;
wire n8673_1;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8678_1;
wire n868;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8683_1;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8688_1;
wire n8689;
wire n8690;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8702;
wire n8702_1;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8707_1;
wire n8709;
wire n8710;
wire n8712;
wire n8712_1;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8717_1;
wire n8718;
wire n8719;
wire n8720;
wire n8721;
wire n8722;
wire n8722_1;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8727_1;
wire n8728;
wire n8729;
wire n873;
wire n8730;
wire n8731;
wire n8732;
wire n8732_1;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8737_1;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8747_1;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8752_1;
wire n8753;
wire n8754;
wire n8756;
wire n8757;
wire n8757_1;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8762_1;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8767_1;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8772_1;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8777_1;
wire n8778;
wire n8779;
wire n878;
wire n8780;
wire n8781;
wire n8782;
wire n8782_1;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8787_1;
wire n8788;
wire n8789;
wire n8790;
wire n8792;
wire n8793;
wire n8794;
wire n8796;
wire n8796_1;
wire n8797;
wire n8799;
wire n8800;
wire n8800_1;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8809;
wire n8809_1;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8814_1;
wire n8815;
wire n8816;
wire n8817;
wire n8819;
wire n8819_1;
wire n8821;
wire n8822;
wire n8824;
wire n8824_1;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8829_1;
wire n883;
wire n8830;
wire n8831;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8839_1;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8844_1;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8852;
wire n8853;
wire n8853_1;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8857_1;
wire n8858;
wire n8859;
wire n8860;
wire n8861;
wire n8862;
wire n8862_1;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8867;
wire n8867_1;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8872_1;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8876_1;
wire n8877;
wire n8878;
wire n8879;
wire n888;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8926;
wire n8929;
wire n893;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8953;
wire n8954;
wire n8955;
wire n8957;
wire n8958;
wire n8959;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8973;
wire n8974;
wire n8975;
wire n8976;
wire n8978;
wire n8979;
wire n898;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8995;
wire n8997;
wire n8998;
wire n8999;
wire n9001;
wire n9002;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9016;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n903;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9058;
wire n9059;
wire n9061;
wire n9062;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9075;
wire n9077;
wire n9078;
wire n9079;
wire n908;
wire n9080;
wire n9081;
wire n9082;
wire n9083;
wire n9084;
wire n9085;
wire n9086;
wire n9087;
wire n9088;
wire n9089;
wire n9090;
wire n9091;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9097;
wire n9098;
wire n9099;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9107;
wire n9108;
wire n9109;
wire n9110;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n913;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9144;
wire n9145;
wire n9146;
wire n9148;
wire n9150;
wire n9151;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9157;
wire n9159;
wire n9160;
wire n9162;
wire n9164;
wire n9165;
wire n9166;
wire n9168;
wire n9169;
wire n917;
wire n9171;
wire n9172;
wire n9173;
wire n9174;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9193;
wire n9194;
wire n9195;
wire n9196;
wire n9197;
wire n9198;
wire n9199;
wire n9200;
wire n9201;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9212;
wire n9213;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9218;
wire n9219;
wire n922;
wire n9220;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9226;
wire n9227;
wire n9229;
wire n9230;
wire n9232;
wire n9234;
wire n9235;
wire n9237;
wire n9238;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9243;
wire n9244;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n9250;
wire n9251;
wire n9253;
wire n9255;
wire n9256;
wire n9257;
wire n9258;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9266;
wire n9267;
wire n9268;
wire n9269;
wire n927;
wire n9270;
wire n9271;
wire n9273;
wire n9274;
wire n9275;
wire n9277;
wire n9278;
wire n9279;
wire n9280;
wire n9281;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9288;
wire n9289;
wire n9290;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9295;
wire n9296;
wire n9297;
wire n9299;
wire n9300;
wire n9301;
wire n9303;
wire n9304;
wire n9306;
wire n9307;
wire n9308;
wire n9310;
wire n9311;
wire n9313;
wire n9314;
wire n9316;
wire n9317;
wire n9318;
wire n9319;
wire n932;
wire n9321;
wire n9322;
wire n9323;
wire n9324;
wire n9325;
wire n9326;
wire n9327;
wire n9328;
wire n9329;
wire n9330;
wire n9331;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9340;
wire n9342;
wire n9343;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9349;
wire n9351;
wire n9352;
wire n9353;
wire n9355;
wire n9357;
wire n9358;
wire n9359;
wire n936;
wire n9360;
wire n9361;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9366;
wire n9367;
wire n9368;
wire n9369;
wire n9371;
wire n9372;
wire n9373;
wire n9374;
wire n9375;
wire n9376;
wire n9377;
wire n9378;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9385;
wire n9387;
wire n9388;
wire n9390;
wire n9392;
wire n9393;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9399;
wire n940;
wire n9400;
wire n9401;
wire n9402;
wire n9403;
wire n9404;
wire n9405;
wire n9406;
wire n9407;
wire n9409;
wire n9410;
wire n9412;
wire n9413;
wire n9414;
wire n9416;
wire n9417;
wire n9418;
wire n9419;
wire n9420;
wire n9421;
wire n9422;
wire n9423;
wire n9425;
wire n9427;
wire n9429;
wire n9431;
wire n9432;
wire n9434;
wire n9435;
wire n9437;
wire n9438;
wire n9439;
wire n9440;
wire n9441;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9447;
wire n9448;
wire n9449;
wire n945;
wire n9450;
wire n9451;
wire n9452;
wire n9454;
wire n9455;
wire n9456;
wire n9457;
wire n9458;
wire n9459;
wire n9460;
wire n9461;
wire n9462;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9468;
wire n9469;
wire n9470;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9476;
wire n9477;
wire n9478;
wire n9480;
wire n9481;
wire n9482;
wire n9484;
wire n9485;
wire n9487;
wire n9488;
wire n9489;
wire n949;
wire n9490;
wire n9491;
wire n9492;
wire n9493;
wire n9494;
wire n9495;
wire n9496;
wire n9497;
wire n9498;
wire n9499;
wire n9500;
wire n9502;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9509;
wire n9510;
wire n9512;
wire n9513;
wire n9514;
wire n9516;
wire n9518;
wire n9520;
wire n9521;
wire n9522;
wire n9523;
wire n9524;
wire n9525;
wire n9526;
wire n9528;
wire n9529;
wire n9531;
wire n9532;
wire n9533;
wire n9535;
wire n9536;
wire n9539;
wire n954;
wire n9540;
wire n9541;
wire n9542;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9547;
wire n9548;
wire n9549;
wire n9550;
wire n9551;
wire n9552;
wire n9553;
wire n9554;
wire n9556;
wire n9557;
wire n9558;
wire n9559;
wire n9560;
wire n9561;
wire n9562;
wire n9563;
wire n9566;
wire n9567;
wire n9568;
wire n9569;
wire n9570;
wire n9571;
wire n9573;
wire n9574;
wire n9575;
wire n9577;
wire n9579;
wire n958;
wire n9580;
wire n9581;
wire n9582;
wire n9584;
wire n9586;
wire n9587;
wire n9588;
wire n9590;
wire n9591;
wire n9592;
wire n9594;
wire n9595;
wire n9597;
wire n9598;
wire n9600;
wire n9601;
wire n9603;
wire n9604;
wire n9606;
wire n9607;
wire n9608;
wire n9609;
wire n9610;
wire n9611;
wire n9612;
wire n9614;
wire n9615;
wire n9617;
wire n9619;
wire n9620;
wire n9621;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9628;
wire n9629;
wire n963;
wire n9630;
wire n9632;
wire n9634;
wire n9635;
wire n9636;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9643;
wire n9644;
wire n9645;
wire n9647;
wire n9648;
wire n9650;
wire n9651;
wire n9652;
wire n9655;
wire n9656;
wire n9657;
wire n9658;
wire n9659;
wire n9660;
wire n9661;
wire n9662;
wire n9663;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9676;
wire n9677;
wire n9678;
wire n9679;
wire n968;
wire n9680;
wire n9681;
wire n9682;
wire n9683;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
wire n9689;
wire n9691;
wire n9693;
wire n9694;
wire n9696;
wire n9698;
wire n9699;
wire n9700;
wire n9701;
wire n9702;
wire n9703;
wire n9704;
wire n9705;
wire n9706;
wire n9707;
wire n9708;
wire n9709;
wire n9710;
wire n9711;
wire n9712;
wire n9713;
wire n9714;
wire n9715;
wire n9716;
wire n9717;
wire n9718;
wire n9719;
wire n9720;
wire n9721;
wire n9722;
wire n9723;
wire n9724;
wire n9725;
wire n9726;
wire n9727;
wire n9728;
wire n9729;
wire n973;
wire n9730;
wire n9731;
wire n9732;
wire n9733;
wire n9734;
wire n9735;
wire n9736;
wire n9738;
wire n9741;
wire n9742;
wire n9745;
wire n9747;
wire n9748;
wire n9750;
wire n9752;
wire n9753;
wire n9755;
wire n9756;
wire n9757;
wire n9758;
wire n9759;
wire n9760;
wire n9761;
wire n9762;
wire n9763;
wire n9764;
wire n9765;
wire n9766;
wire n9767;
wire n9768;
wire n9769;
wire n9770;
wire n9771;
wire n9772;
wire n9773;
wire n9774;
wire n9775;
wire n9776;
wire n9777;
wire n9779;
wire n978;
wire n9780;
wire n9781;
wire n9782;
wire n9784;
wire n9786;
wire n9787;
wire n9788;
wire n9789;
wire n9790;
wire n9791;
wire n9792;
wire n9793;
wire n9794;
wire n9795;
wire n9796;
wire n9798;
wire n9799;
wire n9800;
wire n9802;
wire n9803;
wire n9804;
wire n9805;
wire n9806;
wire n9807;
wire n9810;
wire n9811;
wire n9812;
wire n9813;
wire n9814;
wire n9815;
wire n9816;
wire n9817;
wire n9818;
wire n9819;
wire n982;
wire n9820;
wire n9821;
wire n9822;
wire n9823;
wire n9825;
wire n9826;
wire n9827;
wire n9828;
wire n9829;
wire n9830;
wire n9831;
wire n9833;
wire n9834;
wire n9835;
wire n9836;
wire n9837;
wire n9838;
wire n9839;
wire n9840;
wire n9841;
wire n9843;
wire n9844;
wire n9845;
wire n9846;
wire n9847;
wire n9848;
wire n9849;
wire n9850;
wire n9851;
wire n9852;
wire n9853;
wire n9854;
wire n9855;
wire n9856;
wire n9857;
wire n9858;
wire n9859;
wire n9860;
wire n9861;
wire n9862;
wire n9863;
wire n9864;
wire n9865;
wire n9866;
wire n9867;
wire n9868;
wire n9869;
wire n987;
wire n9870;
wire n9871;
wire n9872;
wire n9873;
wire n9874;
wire n9875;
wire n9876;
wire n9877;
wire n9878;
wire n9879;
wire n9880;
wire n9881;
wire n9882;
wire n9883;
wire n9884;
wire n9887;
wire n9888;
wire n9889;
wire n9891;
wire n9893;
wire n9894;
wire n9895;
wire n9897;
wire n9898;
wire n9900;
wire n9901;
wire n9903;
wire n9904;
wire n9905;
wire n9906;
wire n9907;
wire n9908;
wire n9909;
wire n9910;
wire n9911;
wire n9912;
wire n9913;
wire n9914;
wire n9915;
wire n9916;
wire n9917;
wire n9918;
wire n9919;
wire n992;
wire n9920;
wire n9922;
wire n9923;
wire n9924;
wire n9926;
wire n9927;
wire n9928;
wire n9929;
wire n9930;
wire n9931;
wire n9932;
wire n9933;
wire n9935;
wire n9936;
wire n9937;
wire n9939;
wire n9940;
wire n9941;
wire n9943;
wire n9944;
wire n9945;
wire n9946;
wire n9947;
wire n9948;
wire n9949;
wire n9950;
wire n9952;
wire n9953;
wire n9954;
wire n9956;
wire n9958;
wire n9960;
wire n9963;
wire n9964;
wire n9965;
wire n9967;
wire n9968;
wire n997;
wire n9970;
wire n9971;
wire n9972;
wire n9974;
wire n9975;
wire n9976;
wire n9977;
wire n9978;
wire n9979;
wire n9980;
wire n9981;
wire n9982;
wire n9983;
wire n9984;
wire n9985;
wire n9986;
wire n9988;
wire n9989;
wire n9991;
wire n9993;
wire n9994;
wire n9995;
wire n9996;
wire n9997;
wire n9998;
wire n9999;
wire net_100;
wire net_10000;
wire net_10001;
wire net_10002;
wire net_10003;
wire net_10004;
wire net_10005;
wire net_10006;
wire net_10007;
wire net_10008;
wire net_10009;
wire net_10010;
wire net_10011;
wire net_10012;
wire net_10013;
wire net_10014;
wire net_10015;
wire net_10016;
wire net_10017;
wire net_10018;
wire net_10019;
wire net_10020;
wire net_10021;
wire net_10022;
wire net_10023;
wire net_10024;
wire net_10034;
wire net_10035;
wire net_10036;
wire net_10038;
wire net_10039;
wire net_10044;
wire net_10045;
wire net_10046;
wire net_10047;
wire net_10050;
wire net_10051;
wire net_10052;
wire net_10053;
wire net_10058;
wire net_10059;
wire net_10060;
wire net_10063;
wire net_10064;
wire net_10065;
wire net_10066;
wire net_10067;
wire net_10068;
wire net_10069;
wire net_10070;
wire net_10071;
wire net_10072;
wire net_10073;
wire net_10074;
wire net_10075;
wire net_10076;
wire net_10077;
wire net_10078;
wire net_10079;
wire net_10080;
wire net_10081;
wire net_10082;
wire net_10083;
wire net_10084;
wire net_10085;
wire net_10086;
wire net_10087;
wire net_10088;
wire net_10089;
wire net_10093;
wire net_101;
wire net_10132;
wire net_10133;
wire net_10134;
wire net_10135;
wire net_10169;
wire net_10170;
wire net_10175;
wire net_10176;
wire net_10177;
wire net_10178;
wire net_10179;
wire net_10180;
wire net_10181;
wire net_10182;
wire net_10183;
wire net_10184;
wire net_10185;
wire net_10186;
wire net_10187;
wire net_10188;
wire net_10189;
wire net_10190;
wire net_10191;
wire net_10192;
wire net_10193;
wire net_10194;
wire net_10195;
wire net_10198;
wire net_10199;
wire net_102;
wire net_10237;
wire net_10238;
wire net_10239;
wire net_10240;
wire net_10274;
wire net_10275;
wire net_10280;
wire net_10281;
wire net_10282;
wire net_10283;
wire net_10284;
wire net_10285;
wire net_10286;
wire net_10287;
wire net_10288;
wire net_10289;
wire net_10290;
wire net_10291;
wire net_10292;
wire net_10293;
wire net_10294;
wire net_10295;
wire net_10296;
wire net_10297;
wire net_10298;
wire net_10299;
wire net_103;
wire net_10300;
wire net_10303;
wire net_10304;
wire net_10342;
wire net_10343;
wire net_10344;
wire net_10345;
wire net_10379;
wire net_10380;
wire net_10385;
wire net_10386;
wire net_10387;
wire net_10388;
wire net_10389;
wire net_10390;
wire net_10391;
wire net_10392;
wire net_10393;
wire net_10394;
wire net_10395;
wire net_10396;
wire net_10397;
wire net_10398;
wire net_10399;
wire net_104;
wire net_10400;
wire net_10401;
wire net_10402;
wire net_10403;
wire net_10404;
wire net_10405;
wire net_10408;
wire net_10409;
wire net_10447;
wire net_10448;
wire net_10449;
wire net_10450;
wire net_10484;
wire net_10485;
wire net_10490;
wire net_10491;
wire net_10492;
wire net_10493;
wire net_10494;
wire net_10495;
wire net_10496;
wire net_10497;
wire net_10498;
wire net_10499;
wire net_105;
wire net_10500;
wire net_10501;
wire net_10502;
wire net_10503;
wire net_10504;
wire net_10505;
wire net_10506;
wire net_10507;
wire net_10508;
wire net_10509;
wire net_10510;
wire net_10513;
wire net_10514;
wire net_10516;
wire net_10517;
wire net_10518;
wire net_10519;
wire net_10520;
wire net_10521;
wire net_10522;
wire net_10523;
wire net_10524;
wire net_10525;
wire net_10526;
wire net_10527;
wire net_10530;
wire net_10532;
wire net_10533;
wire net_10536;
wire net_10537;
wire net_10539;
wire net_10540;
wire net_10541;
wire net_10542;
wire net_106;
wire net_107;
wire net_108;
wire net_109;
wire net_110;
wire net_111;
wire net_112;
wire net_113;
wire net_114;
wire net_115;
wire net_116;
wire net_134;
wire net_135;
wire net_136;
wire net_137;
wire net_138;
wire net_139;
wire net_140;
wire net_141;
wire net_142;
wire net_143;
wire net_144;
wire net_145;
wire net_146;
wire net_147;
wire net_148;
wire net_149;
wire net_150;
wire net_186;
wire net_192;
wire net_194;
wire net_195;
wire net_196;
wire net_197;
wire net_203;
wire net_204;
wire net_205;
wire net_206;
wire net_207;
wire net_208;
wire net_209;
wire net_210;
wire net_211;
wire net_212;
wire net_213;
wire net_214;
wire net_215;
wire net_216;
wire net_217;
wire net_218;
wire net_219;
wire net_220;
wire net_221;
wire net_222;
wire net_223;
wire net_224;
wire net_225;
wire net_226;
wire net_227;
wire net_228;
wire net_229;
wire net_230;
wire net_235;
wire net_236;
wire net_237;
wire net_238;
wire net_239;
wire net_240;
wire net_241;
wire net_242;
wire net_243;
wire net_244;
wire net_245;
wire net_246;
wire net_247;
wire net_248;
wire net_249;
wire net_250;
wire net_251;
wire net_252;
wire net_253;
wire net_256;
wire net_257;
wire net_258;
wire net_260;
wire net_262;
wire net_263;
wire net_264;
wire net_279;
wire net_281;
wire net_282;
wire net_283;
wire net_284;
wire net_285;
wire net_286;
wire net_287;
wire net_288;
wire net_289;
wire net_290;
wire net_291;
wire net_292;
wire net_293;
wire net_294;
wire net_295;
wire net_296;
wire net_297;
wire net_298;
wire net_299;
wire net_300;
wire net_301;
wire net_302;
wire net_303;
wire net_304;
wire net_305;
wire net_306;
wire net_307;
wire net_308;
wire net_309;
wire net_310;
wire net_311;
wire net_312;
wire net_313;
wire net_8816;
wire net_8818;
wire net_8820;
wire net_8822;
wire net_8827;
wire net_8832;
wire net_8835;
wire net_8836;
wire net_8837;
wire net_8838;
wire net_90;
wire net_91;
wire net_9116;
wire net_9119;
wire net_9120;
wire net_9121;
wire net_9122;
wire net_9123;
wire net_9124;
wire net_9125;
wire net_9126;
wire net_9127;
wire net_9128;
wire net_9129;
wire net_9130;
wire net_9131;
wire net_9132;
wire net_9133;
wire net_9134;
wire net_9135;
wire net_9136;
wire net_9137;
wire net_9138;
wire net_9139;
wire net_9140;
wire net_9141;
wire net_9142;
wire net_9143;
wire net_9144;
wire net_9145;
wire net_9146;
wire net_9147;
wire net_9148;
wire net_9149;
wire net_9150;
wire net_9151;
wire net_9152;
wire net_9153;
wire net_9154;
wire net_9155;
wire net_9156;
wire net_9157;
wire net_9158;
wire net_9159;
wire net_9162;
wire net_9163;
wire net_9170;
wire net_9174;
wire net_9175;
wire net_9179;
wire net_9180;
wire net_9181;
wire net_9182;
wire net_9184;
wire net_9197;
wire net_9198;
wire net_9199;
wire net_92;
wire net_9200;
wire net_9205;
wire net_9206;
wire net_9208;
wire net_9210;
wire net_9212;
wire net_9216;
wire net_9218;
wire net_9219;
wire net_9220;
wire net_9221;
wire net_9222;
wire net_9223;
wire net_9224;
wire net_9225;
wire net_9226;
wire net_9227;
wire net_9228;
wire net_9229;
wire net_9230;
wire net_9231;
wire net_9233;
wire net_9234;
wire net_9251;
wire net_9252;
wire net_9253;
wire net_9254;
wire net_9255;
wire net_9256;
wire net_9257;
wire net_9259;
wire net_9260;
wire net_9261;
wire net_9262;
wire net_9263;
wire net_9264;
wire net_9265;
wire net_9269;
wire net_9270;
wire net_9271;
wire net_9273;
wire net_9274;
wire net_9275;
wire net_9276;
wire net_9277;
wire net_9278;
wire net_9279;
wire net_9280;
wire net_9281;
wire net_9282;
wire net_9283;
wire net_9284;
wire net_9285;
wire net_9286;
wire net_9287;
wire net_9288;
wire net_9289;
wire net_93;
wire net_9303;
wire net_9304;
wire net_9305;
wire net_9306;
wire net_9307;
wire net_9308;
wire net_9310;
wire net_9327;
wire net_9328;
wire net_9329;
wire net_9330;
wire net_9331;
wire net_9332;
wire net_9333;
wire net_9334;
wire net_9335;
wire net_9336;
wire net_9337;
wire net_9338;
wire net_9339;
wire net_9340;
wire net_9341;
wire net_9342;
wire net_9347;
wire net_9348;
wire net_9349;
wire net_9350;
wire net_9357;
wire net_9358;
wire net_9359;
wire net_9360;
wire net_9361;
wire net_9364;
wire net_9365;
wire net_9366;
wire net_9367;
wire net_9368;
wire net_9369;
wire net_9379;
wire net_9387;
wire net_94;
wire net_9425;
wire net_9426;
wire net_9430;
wire net_9431;
wire net_9432;
wire net_9433;
wire net_9435;
wire net_9436;
wire net_9438;
wire net_9439;
wire net_9440;
wire net_9441;
wire net_9442;
wire net_9443;
wire net_9444;
wire net_9445;
wire net_9446;
wire net_9447;
wire net_9448;
wire net_9449;
wire net_9450;
wire net_9451;
wire net_9452;
wire net_9453;
wire net_9454;
wire net_9455;
wire net_9456;
wire net_9457;
wire net_9458;
wire net_9459;
wire net_9460;
wire net_9461;
wire net_9462;
wire net_9463;
wire net_9464;
wire net_9465;
wire net_9466;
wire net_9467;
wire net_9468;
wire net_9469;
wire net_9470;
wire net_9471;
wire net_9472;
wire net_9473;
wire net_9474;
wire net_9475;
wire net_9476;
wire net_9477;
wire net_9478;
wire net_9479;
wire net_9480;
wire net_9481;
wire net_9482;
wire net_9483;
wire net_9484;
wire net_9485;
wire net_9486;
wire net_9487;
wire net_9488;
wire net_9489;
wire net_9490;
wire net_9491;
wire net_9492;
wire net_9493;
wire net_9494;
wire net_9495;
wire net_9496;
wire net_9497;
wire net_9498;
wire net_9499;
wire net_95;
wire net_9500;
wire net_9501;
wire net_9504;
wire net_9505;
wire net_9506;
wire net_9507;
wire net_9508;
wire net_9509;
wire net_9510;
wire net_9511;
wire net_9513;
wire net_9522;
wire net_9523;
wire net_9524;
wire net_9525;
wire net_9526;
wire net_9527;
wire net_9528;
wire net_9529;
wire net_9531;
wire net_9533;
wire net_9534;
wire net_9535;
wire net_9538;
wire net_9539;
wire net_9540;
wire net_9542;
wire net_9543;
wire net_9544;
wire net_9545;
wire net_9549;
wire net_9559;
wire net_9560;
wire net_9568;
wire net_9570;
wire net_9571;
wire net_9574;
wire net_9575;
wire net_9576;
wire net_9577;
wire net_9578;
wire net_9579;
wire net_9582;
wire net_9583;
wire net_9584;
wire net_9585;
wire net_9586;
wire net_9587;
wire net_9592;
wire net_9593;
wire net_9594;
wire net_9595;
wire net_9596;
wire net_9597;
wire net_9598;
wire net_9599;
wire net_96;
wire net_9604;
wire net_9605;
wire net_9607;
wire net_9610;
wire net_9612;
wire net_9613;
wire net_9614;
wire net_9615;
wire net_9616;
wire net_9617;
wire net_9618;
wire net_9619;
wire net_9620;
wire net_9621;
wire net_9622;
wire net_9623;
wire net_9624;
wire net_9625;
wire net_9626;
wire net_9631;
wire net_9632;
wire net_9634;
wire net_9647;
wire net_9648;
wire net_9650;
wire net_9651;
wire net_9652;
wire net_9653;
wire net_9654;
wire net_9655;
wire net_9656;
wire net_9657;
wire net_9659;
wire net_9662;
wire net_9663;
wire net_9664;
wire net_9665;
wire net_9666;
wire net_9667;
wire net_9668;
wire net_9669;
wire net_9670;
wire net_9671;
wire net_9672;
wire net_9673;
wire net_9674;
wire net_9675;
wire net_9676;
wire net_9677;
wire net_9678;
wire net_9679;
wire net_9680;
wire net_9681;
wire net_9682;
wire net_9683;
wire net_9684;
wire net_9685;
wire net_9686;
wire net_9687;
wire net_9688;
wire net_9689;
wire net_9690;
wire net_9691;
wire net_9692;
wire net_9693;
wire net_9694;
wire net_9695;
wire net_9696;
wire net_9697;
wire net_9698;
wire net_9699;
wire net_97;
wire net_9700;
wire net_9701;
wire net_9702;
wire net_9703;
wire net_9704;
wire net_9705;
wire net_9706;
wire net_9707;
wire net_9708;
wire net_9709;
wire net_9710;
wire net_9711;
wire net_9712;
wire net_9713;
wire net_9714;
wire net_9715;
wire net_9716;
wire net_9717;
wire net_9718;
wire net_9719;
wire net_9720;
wire net_9721;
wire net_9722;
wire net_9723;
wire net_9724;
wire net_9725;
wire net_9726;
wire net_9727;
wire net_9737;
wire net_9738;
wire net_9739;
wire net_9741;
wire net_9742;
wire net_9747;
wire net_9748;
wire net_9749;
wire net_9750;
wire net_9753;
wire net_9754;
wire net_9755;
wire net_9756;
wire net_9757;
wire net_9758;
wire net_9759;
wire net_9760;
wire net_9761;
wire net_9762;
wire net_9763;
wire net_9764;
wire net_9765;
wire net_9766;
wire net_9767;
wire net_9768;
wire net_9769;
wire net_9770;
wire net_9771;
wire net_9772;
wire net_9773;
wire net_9774;
wire net_9775;
wire net_9776;
wire net_9777;
wire net_9778;
wire net_9779;
wire net_9780;
wire net_9781;
wire net_9782;
wire net_9783;
wire net_9784;
wire net_9785;
wire net_9786;
wire net_9787;
wire net_9788;
wire net_9789;
wire net_9790;
wire net_9791;
wire net_9792;
wire net_9793;
wire net_9794;
wire net_9795;
wire net_9796;
wire net_9797;
wire net_9798;
wire net_9799;
wire net_98;
wire net_9800;
wire net_9801;
wire net_9802;
wire net_9803;
wire net_9804;
wire net_9805;
wire net_9806;
wire net_9807;
wire net_9808;
wire net_9809;
wire net_9810;
wire net_9811;
wire net_9812;
wire net_9813;
wire net_9814;
wire net_9815;
wire net_9816;
wire net_9817;
wire net_9818;
wire net_9819;
wire net_9820;
wire net_9821;
wire net_9822;
wire net_9823;
wire net_9824;
wire net_9825;
wire net_9826;
wire net_9836;
wire net_9837;
wire net_9838;
wire net_9840;
wire net_9841;
wire net_9846;
wire net_9847;
wire net_9848;
wire net_9849;
wire net_9852;
wire net_9853;
wire net_9854;
wire net_9855;
wire net_9856;
wire net_9857;
wire net_9858;
wire net_9859;
wire net_9860;
wire net_9861;
wire net_9862;
wire net_9863;
wire net_9864;
wire net_9865;
wire net_9866;
wire net_9867;
wire net_9868;
wire net_9869;
wire net_9870;
wire net_9871;
wire net_9872;
wire net_9873;
wire net_9874;
wire net_9875;
wire net_9876;
wire net_9877;
wire net_9878;
wire net_9879;
wire net_9880;
wire net_9881;
wire net_9882;
wire net_9883;
wire net_9884;
wire net_9885;
wire net_9886;
wire net_9887;
wire net_9888;
wire net_9889;
wire net_9890;
wire net_9891;
wire net_9892;
wire net_9893;
wire net_9894;
wire net_9895;
wire net_9896;
wire net_9897;
wire net_9898;
wire net_9899;
wire net_99;
wire net_9900;
wire net_9901;
wire net_9902;
wire net_9903;
wire net_9904;
wire net_9905;
wire net_9906;
wire net_9907;
wire net_9908;
wire net_9909;
wire net_9910;
wire net_9911;
wire net_9912;
wire net_9913;
wire net_9914;
wire net_9915;
wire net_9916;
wire net_9917;
wire net_9918;
wire net_9919;
wire net_9920;
wire net_9921;
wire net_9922;
wire net_9923;
wire net_9924;
wire net_9925;
wire net_9935;
wire net_9936;
wire net_9937;
wire net_9939;
wire net_9940;
wire net_9945;
wire net_9946;
wire net_9947;
wire net_9948;
wire net_9951;
wire net_9952;
wire net_9953;
wire net_9954;
wire net_9955;
wire net_9956;
wire net_9959;
wire net_9960;
wire net_9961;
wire net_9962;
wire net_9963;
wire net_9964;
wire net_9965;
wire net_9966;
wire net_9967;
wire net_9968;
wire net_9969;
wire net_9970;
wire net_9971;
wire net_9972;
wire net_9973;
wire net_9974;
wire net_9975;
wire net_9976;
wire net_9977;
wire net_9978;
wire net_9979;
wire net_9980;
wire net_9981;
wire net_9982;
wire net_9983;
wire net_9984;
wire net_9985;
wire net_9986;
wire net_9987;
wire net_9988;
wire net_9989;
wire net_9990;
wire net_9991;
wire net_9992;
wire net_9993;
wire net_9994;
wire net_9995;
wire net_9996;
wire net_9997;
wire net_9998;
wire net_9999;
wire x185128;
wire x185129;
wire x185130;
wire x185131;
wire x185132;
wire x185133;
wire x185134;
wire x185135;
wire x185136;
wire x185137;
wire x185138;
wire x185139;
wire x185140;
wire x185141;
wire x3675;

// Start cells
in01f01  g0000 ( .o(n5488), .a(x4587) );
in01f01  g0001 ( .o(n5489), .a(_net_9437) );
na02f01  g0002 ( .o(n5490), .a(_net_9532), .b(n5489) );
no02f01  g0003 ( .o(n7916), .a(n5490), .b(_net_9250) );
no03f01  g0004 ( .o(n5492), .a(n7916), .b(_net_9537), .c(_net_9536) );
no02f01  g0005 ( .o(n5493), .a(n5492), .b(_net_9437) );
no02f01  g0006 ( .o(n5494), .a(n5493), .b(_net_9541) );
in01f01  g0007 ( .o(n5495_1), .a(_net_10529) );
na02f01  g0008 ( .o(n5496), .a(n5494), .b(_net_9658) );
in01f01  g0009 ( .o(n5497), .a(n5496) );
no02f01  g0010 ( .o(n5498), .a(_net_10531), .b(net_10530) );
in01f01  g0011 ( .o(n5499), .a(x6157) );
in01f01  g0012 ( .o(n5500_1), .a(x3867) );
in01f01  g0013 ( .o(n5501), .a(_net_10538) );
no03f01  g0014 ( .o(n5502), .a(n5501), .b(n5500_1), .c(n5499) );
no03f01  g0015 ( .o(n5503), .a(n5501), .b(x3867), .c(n5499) );
no02f01  g0016 ( .o(n5504_1), .a(n5503), .b(n5502) );
oa22f01  g0017 ( .o(n5505), .a(n5504_1), .b(n5495_1), .c(n5498), .d(n5497) );
oa12f01  g0018 ( .o(n5506), .a(n5494), .b(n5505), .c(_net_9658) );
na02f01  g0019 ( .o(n5507), .a(n5506), .b(net_303) );
oa12f01  g0020 ( .o(x91), .a(n5507), .b(n5506), .c(n5488) );
in01f01  g0021 ( .o(n5509), .a(_net_277) );
in01f01  g0022 ( .o(n5510), .a(n5506) );
na02f01  g0023 ( .o(n5511), .a(n5510), .b(x6220) );
oa12f01  g0024 ( .o(x329), .a(n5511), .b(n5510), .c(n5509) );
in01f01  g0025 ( .o(n5513_1), .a(x6028) );
na02f01  g0026 ( .o(n5514), .a(n5506), .b(net_282) );
oa12f01  g0027 ( .o(x293), .a(n5514), .b(n5506), .c(n5513_1) );
in01f01  g0028 ( .o(n5516), .a(x4520) );
na02f01  g0029 ( .o(n5517), .a(n5506), .b(net_304) );
oa12f01  g0030 ( .o(x86), .a(n5517), .b(n5506), .c(n5516) );
in01f01  g0031 ( .o(n5519), .a(x3507) );
in01f01  g0032 ( .o(n5520), .a(_net_10543) );
oa22f01  g0033 ( .o(x507), .a(net_9233), .b(n5520), .c(n5519), .d(x3534) );
in01f01  g0034 ( .o(n5522), .a(_net_274) );
na02f01  g0035 ( .o(n5523_1), .a(n5510), .b(x6264) );
oa12f01  g0036 ( .o(x355), .a(n5523_1), .b(n5510), .c(n5522) );
in01f01  g0037 ( .o(n5525), .a(x4041) );
na02f01  g0038 ( .o(n5526), .a(n5506), .b(net_310) );
oa12f01  g0039 ( .o(x39), .a(n5526), .b(n5506), .c(n5525) );
in01f01  g0040 ( .o(n5528_1), .a(_net_271) );
na02f01  g0041 ( .o(n5529), .a(n5510), .b(x6327) );
oa12f01  g0042 ( .o(x381), .a(n5529), .b(n5510), .c(n5528_1) );
in01f01  g0043 ( .o(n5531), .a(x5225) );
na02f01  g0044 ( .o(n5532), .a(n5506), .b(net_295) );
oa12f01  g0045 ( .o(x143), .a(n5532), .b(n5506), .c(n5531) );
in01f01  g0046 ( .o(n5534), .a(_net_275) );
na02f01  g0047 ( .o(n5535), .a(n5510), .b(x6252) );
oa12f01  g0048 ( .o(x348), .a(n5535), .b(n5510), .c(n5534) );
in01f01  g0049 ( .o(n5537_1), .a(x5790) );
na02f01  g0050 ( .o(n5538), .a(n5506), .b(net_286) );
oa12f01  g0051 ( .o(x257), .a(n5538), .b(n5506), .c(n5537_1) );
in01f01  g0052 ( .o(n5540), .a(x5901) );
na02f01  g0053 ( .o(n5541), .a(n5506), .b(net_284) );
oa12f01  g0054 ( .o(x277), .a(n5541), .b(n5506), .c(n5540) );
in01f01  g0055 ( .o(n5543), .a(_net_278) );
na02f01  g0056 ( .o(n5544), .a(n5510), .b(x6198) );
oa12f01  g0057 ( .o(x316), .a(n5544), .b(n5510), .c(n5543) );
in01f01  g0058 ( .o(n5546), .a(x4851) );
na02f01  g0059 ( .o(n5547_1), .a(n5506), .b(net_300) );
oa12f01  g0060 ( .o(x111), .a(n5547_1), .b(n5506), .c(n5546) );
in01f01  g0061 ( .o(n5549), .a(x6496) );
na02f01  g0062 ( .o(n5550), .a(n5506), .b(_net_267) );
oa12f01  g0063 ( .o(x420), .a(n5550), .b(n5506), .c(n5549) );
in01f01  g0064 ( .o(n5552_1), .a(x4694) );
na02f01  g0065 ( .o(n5553), .a(n5506), .b(net_302) );
oa12f01  g0066 ( .o(x101), .a(n5553), .b(n5506), .c(n5552_1) );
in01f01  g0067 ( .o(n5555), .a(x3949) );
na02f01  g0068 ( .o(n5556), .a(n5506), .b(net_311) );
oa12f01  g0069 ( .o(x33), .a(n5556), .b(n5506), .c(n5555) );
in01f01  g0070 ( .o(n5558), .a(x6531) );
na02f01  g0071 ( .o(n5559), .a(n5506), .b(_net_266) );
oa12f01  g0072 ( .o(x427), .a(n5559), .b(n5506), .c(n5558) );
in01f01  g0073 ( .o(n5561), .a(x5722) );
na02f01  g0074 ( .o(n5562_1), .a(n5506), .b(net_287) );
oa12f01  g0075 ( .o(x244), .a(n5562_1), .b(n5506), .c(n5561) );
in01f01  g0076 ( .o(n5564), .a(x6401) );
na02f01  g0077 ( .o(n5565), .a(n5506), .b(_net_269) );
oa12f01  g0078 ( .o(x401), .a(n5565), .b(n5506), .c(n5564) );
in01f01  g0079 ( .o(n5567_1), .a(x4359) );
na02f01  g0080 ( .o(n5568), .a(n5506), .b(net_306) );
oa12f01  g0081 ( .o(x73), .a(n5568), .b(n5506), .c(n5567_1) );
in01f01  g0082 ( .o(n5570), .a(x6102) );
na02f01  g0083 ( .o(n5571), .a(n5506), .b(net_281) );
oa12f01  g0084 ( .o(x297), .a(n5571), .b(n5506), .c(n5570) );
in01f01  g0085 ( .o(n5573), .a(x5850) );
na02f01  g0086 ( .o(n5574), .a(n5506), .b(net_285) );
oa12f01  g0087 ( .o(x268), .a(n5574), .b(n5506), .c(n5573) );
in01f01  g0088 ( .o(n5576), .a(x5077) );
na02f01  g0089 ( .o(n5577_1), .a(n5506), .b(net_297) );
oa12f01  g0090 ( .o(x126), .a(n5577_1), .b(n5506), .c(n5576) );
in01f01  g0091 ( .o(n5579), .a(_net_276) );
na02f01  g0092 ( .o(n5580), .a(n5510), .b(x6241) );
oa12f01  g0093 ( .o(x341), .a(n5580), .b(n5510), .c(n5579) );
in01f01  g0094 ( .o(n5582_1), .a(x5143) );
na02f01  g0095 ( .o(n5583), .a(n5506), .b(net_296) );
oa12f01  g0096 ( .o(x132), .a(n5583), .b(n5506), .c(n5582_1) );
in01f01  g0097 ( .o(n5585_1), .a(x5498) );
na02f01  g0098 ( .o(n5586), .a(n5506), .b(net_291) );
oa12f01  g0099 ( .o(x198), .a(n5586), .b(n5506), .c(n5585_1) );
in01f01  g0100 ( .o(n5588), .a(_net_272) );
na02f01  g0101 ( .o(n5589_1), .a(n5510), .b(x6303) );
oa12f01  g0102 ( .o(x374), .a(n5589_1), .b(n5510), .c(n5588) );
in01f01  g0103 ( .o(n5591), .a(x5003) );
na02f01  g0104 ( .o(n5592), .a(n5506), .b(net_298) );
oa12f01  g0105 ( .o(x121), .a(n5592), .b(n5506), .c(n5591) );
in01f01  g0106 ( .o(n5594_1), .a(net_279) );
na02f01  g0107 ( .o(n5595), .a(n5510), .b(x6186) );
oa12f01  g0108 ( .o(x304), .a(n5595), .b(n5510), .c(n5594_1) );
in01f01  g0109 ( .o(n5597_1), .a(x4449) );
na02f01  g0110 ( .o(n5598), .a(n5506), .b(net_305) );
oa12f01  g0111 ( .o(x80), .a(n5598), .b(n5506), .c(n5597_1) );
in01f01  g0112 ( .o(n5600), .a(x5427) );
na02f01  g0113 ( .o(n5601_1), .a(n5506), .b(net_292) );
oa12f01  g0114 ( .o(x182), .a(n5601_1), .b(n5506), .c(n5600) );
in01f01  g0115 ( .o(n5603), .a(x5289) );
na02f01  g0116 ( .o(n5604), .a(n5506), .b(net_294) );
oa12f01  g0117 ( .o(x157), .a(n5604), .b(n5506), .c(n5603) );
in01f01  g0118 ( .o(n5606), .a(x5601) );
na02f01  g0119 ( .o(n5607), .a(n5506), .b(net_289) );
oa12f01  g0120 ( .o(x223), .a(n5607), .b(n5506), .c(n5606) );
in01f01  g0121 ( .o(n5609), .a(x4285) );
na02f01  g0122 ( .o(n5610_1), .a(n5506), .b(net_307) );
oa12f01  g0123 ( .o(x65), .a(n5610_1), .b(n5506), .c(n5609) );
in01f01  g0124 ( .o(n5612), .a(x4937) );
na02f01  g0125 ( .o(n5613), .a(n5506), .b(net_299) );
oa12f01  g0126 ( .o(x116), .a(n5613), .b(n5506), .c(n5612) );
in01f01  g0127 ( .o(n5615), .a(x4117) );
na02f01  g0128 ( .o(n5616), .a(n5506), .b(net_309) );
oa12f01  g0129 ( .o(x46), .a(n5616), .b(n5506), .c(n5615) );
in01f01  g0130 ( .o(n5618), .a(x5647) );
na02f01  g0131 ( .o(n5619_1), .a(n5506), .b(net_288) );
oa12f01  g0132 ( .o(x233), .a(n5619_1), .b(n5506), .c(n5618) );
in01f01  g0133 ( .o(n5621), .a(x5961) );
na02f01  g0134 ( .o(n5622), .a(n5506), .b(net_283) );
oa12f01  g0135 ( .o(x285), .a(n5622), .b(n5506), .c(n5621) );
in01f01  g0136 ( .o(n2227), .a(n5494) );
na03f01  g0137 ( .o(n5625), .a(n5506), .b(n2227), .c(_net_314) );
na02f01  g0138 ( .o(n5626), .a(n5496), .b(net_10530) );
na02f01  g0139 ( .o(n5627), .a(n5502), .b(_net_10529) );
na02f01  g0140 ( .o(n5628), .a(n5627), .b(n5626) );
na02f01  g0141 ( .o(n5629_1), .a(n5628), .b(n5505) );
oa12f01  g0142 ( .o(x0), .a(n5625), .b(n5629_1), .c(n5506) );
in01f01  g0143 ( .o(n5631), .a(x6445) );
na02f01  g0144 ( .o(n5632), .a(n5506), .b(_net_268) );
oa12f01  g0145 ( .o(x413), .a(n5632), .b(n5506), .c(n5631) );
in01f01  g0146 ( .o(n5634), .a(x5364) );
na02f01  g0147 ( .o(n5635), .a(n5506), .b(net_293) );
oa12f01  g0148 ( .o(x166), .a(n5635), .b(n5506), .c(n5634) );
in01f01  g0149 ( .o(n5637), .a(x4209) );
na02f01  g0150 ( .o(n5638_1), .a(n5506), .b(net_308) );
oa12f01  g0151 ( .o(x57), .a(n5638_1), .b(n5506), .c(n5637) );
in01f01  g0152 ( .o(n5640), .a(x4781) );
na02f01  g0153 ( .o(n5641), .a(n5506), .b(net_301) );
oa12f01  g0154 ( .o(x106), .a(n5641), .b(n5506), .c(n5640) );
in01f01  g0155 ( .o(n5643), .a(_net_273) );
na02f01  g0156 ( .o(n5644), .a(n5510), .b(x6282) );
oa12f01  g0157 ( .o(x366), .a(n5644), .b(n5510), .c(n5643) );
in01f01  g0158 ( .o(n5646), .a(x3889) );
na02f01  g0159 ( .o(n5647_1), .a(n5506), .b(net_312) );
oa12f01  g0160 ( .o(x27), .a(n5647_1), .b(n5506), .c(n5646) );
in01f01  g0161 ( .o(n5649), .a(x5548) );
na02f01  g0162 ( .o(n5650), .a(n5506), .b(net_290) );
oa12f01  g0163 ( .o(x208), .a(n5650), .b(n5506), .c(n5649) );
in01f01  g0164 ( .o(n5652), .a(_net_270) );
na02f01  g0165 ( .o(n5653), .a(n5510), .b(x6351) );
oa12f01  g0166 ( .o(x389), .a(n5653), .b(n5510), .c(n5652) );
in01f01  g0167 ( .o(n5655), .a(x6577) );
na02f01  g0168 ( .o(n5656_1), .a(n5506), .b(_net_265) );
oa12f01  g0169 ( .o(x437), .a(n5656_1), .b(n5506), .c(n5655) );
in01f01  g0170 ( .o(n5658), .a(x6599) );
no02f01  g0171 ( .o(n5659), .a(n5558), .b(n5655) );
in01f01  g0172 ( .o(n5660), .a(n5659) );
no03f01  g0173 ( .o(n5661_1), .a(n5501), .b(n5500_1), .c(x6157) );
in01f01  g0174 ( .o(n5662), .a(n5661_1) );
no02f01  g0175 ( .o(n5663), .a(n5662), .b(n5495_1) );
in01f01  g0176 ( .o(n5664), .a(n5663) );
no02f01  g0177 ( .o(n5665), .a(x6351), .b(x6327) );
in01f01  g0178 ( .o(n5666_1), .a(n5665) );
no03f01  g0179 ( .o(n5667), .a(n5666_1), .b(x6496), .c(n5564) );
in01f01  g0180 ( .o(n5668), .a(n5667) );
no02f01  g0181 ( .o(n5669), .a(n5668), .b(x6445) );
in01f01  g0182 ( .o(n5670), .a(n5669) );
no02f01  g0183 ( .o(n5671_1), .a(n5670), .b(n5664) );
in01f01  g0184 ( .o(n5672), .a(n5671_1) );
no02f01  g0185 ( .o(n5673), .a(n5672), .b(n5660) );
in01f01  g0186 ( .o(n5674), .a(net_10175) );
no02f01  g0187 ( .o(n5675), .a(_net_9117), .b(_net_166) );
no02f01  g0188 ( .o(n5676_1), .a(n5675), .b(n5674) );
in01f01  g0189 ( .o(n5677), .a(n5676_1) );
no03f01  g0190 ( .o(n5678), .a(n5677), .b(n5673), .c(n5658) );
ao12f01  g0191 ( .o(n5679), .a(n5658), .b(n5678), .c(net_252) );
no03f01  g0192 ( .o(n5680), .a(n5676_1), .b(n5673), .c(n5658) );
no03f01  g0193 ( .o(n5681_1), .a(n5672), .b(n5660), .c(n5658) );
ao22f01  g0194 ( .o(n5682), .a(n5681_1), .b(x4694), .c(n5680), .d(net_9715) );
na02f01  g0195 ( .o(n500), .a(n5682), .b(n5679) );
in01f01  g0196 ( .o(n5684), .a(net_9939) );
no02f01  g0197 ( .o(n5685_1), .a(x6531), .b(x6577) );
in01f01  g0198 ( .o(n5686), .a(n5685_1) );
no02f01  g0199 ( .o(n5687), .a(n5668), .b(n5631) );
in01f01  g0200 ( .o(n5688), .a(n5687) );
no02f01  g0201 ( .o(n5689), .a(n5688), .b(n5664) );
in01f01  g0202 ( .o(n5690_1), .a(n5689) );
no02f01  g0203 ( .o(n5691), .a(n5690_1), .b(n5686) );
na02f01  g0204 ( .o(n5692), .a(n5691), .b(x6599) );
in01f01  g0205 ( .o(n5693), .a(n5691) );
na02f01  g0206 ( .o(n5694), .a(n5693), .b(x6599) );
oa22f01  g0207 ( .o(n505), .a(n5694), .b(n5684), .c(n5692), .d(n5576) );
in01f01  g0208 ( .o(n5696), .a(net_9507) );
in01f01  g0209 ( .o(n5697), .a(_net_9421) );
in01f01  g0210 ( .o(n5698), .a(_net_9062) );
no02f01  g0211 ( .o(n5699), .a(_net_8955), .b(n5698) );
na03f01  g0212 ( .o(n5700_1), .a(n5699), .b(n5697), .c(_net_9512) );
ao12f01  g0213 ( .o(n5701), .a(_net_9421), .b(n5699), .c(_net_9512) );
no02f01  g0214 ( .o(n5702), .a(n5701), .b(n5697) );
ao22f01  g0215 ( .o(n5703), .a(n5702), .b(x2589), .c(n5701), .d(_net_9400) );
oa12f01  g0216 ( .o(n514), .a(n5703), .b(n5700_1), .c(n5696) );
in01f01  g0217 ( .o(n5705_1), .a(_net_9934) );
in01f01  g0218 ( .o(n5706), .a(_net_9927) );
in01f01  g0219 ( .o(n5707), .a(_net_9926) );
oa22f01  g0220 ( .o(n5708), .a(_net_8842), .b(n5707), .c(n5706), .d(_net_10374) );
na02f01  g0221 ( .o(n5709), .a(n5706), .b(_net_10374) );
in01f01  g0222 ( .o(n5710_1), .a(_net_9929) );
in01f01  g0223 ( .o(n5711), .a(_net_9928) );
oa22f01  g0224 ( .o(n5712), .a(_net_10376), .b(n5710_1), .c(n5711), .d(_net_10375) );
ao12f01  g0225 ( .o(n5713), .a(n5712), .b(n5709), .c(n5708) );
in01f01  g0226 ( .o(n5714_1), .a(_net_10376) );
oa12f01  g0227 ( .o(n5715), .a(_net_10375), .b(_net_10376), .c(n5710_1) );
oa22f01  g0228 ( .o(n5716), .a(n5715), .b(_net_9928), .c(n5714_1), .d(_net_9929) );
no02f01  g0229 ( .o(n5717), .a(n5716), .b(n5713) );
in01f01  g0230 ( .o(n5718), .a(_net_9932) );
in01f01  g0231 ( .o(n5719_1), .a(_net_9933) );
oa22f01  g0232 ( .o(n5720), .a(net_10379), .b(n5718), .c(n5719_1), .d(net_10380) );
in01f01  g0233 ( .o(n5721), .a(_net_9930) );
in01f01  g0234 ( .o(n5722), .a(_net_9931) );
oa22f01  g0235 ( .o(n5723), .a(n5722), .b(_net_10378), .c(_net_10377), .d(n5721) );
no03f01  g0236 ( .o(n5724_1), .a(n5723), .b(n5720), .c(n5717) );
in01f01  g0237 ( .o(n5725), .a(_net_10378) );
in01f01  g0238 ( .o(n5726), .a(_net_10377) );
ao12f01  g0239 ( .o(n5727), .a(n5726), .b(_net_9931), .c(n5725) );
ao22f01  g0240 ( .o(n5728), .a(n5727), .b(n5721), .c(n5722), .d(_net_10378) );
oa12f01  g0241 ( .o(n5729_1), .a(net_10379), .b(n5719_1), .c(net_10380) );
no02f01  g0242 ( .o(n5730), .a(n5729_1), .b(_net_9932) );
ao12f01  g0243 ( .o(n5731), .a(n5730), .b(n5719_1), .c(net_10380) );
oa12f01  g0244 ( .o(n5732), .a(n5731), .b(n5728), .c(n5720) );
oa22f01  g0245 ( .o(n5733), .a(n5732), .b(n5724_1), .c(_net_10381), .d(n5705_1) );
na02f01  g0246 ( .o(n5734_1), .a(_net_10381), .b(n5705_1) );
no03f01  g0247 ( .o(n5735), .a(_net_8823), .b(net_8836), .c(net_8822) );
na03f01  g0248 ( .o(n519), .a(n5735), .b(n5734_1), .c(n5733) );
in01f01  g0249 ( .o(n5737), .a(net_9505) );
in01f01  g0250 ( .o(n5738), .a(_net_9512) );
na02f01  g0251 ( .o(n5739_1), .a(_net_8955), .b(_net_9062) );
no02f01  g0252 ( .o(n5740), .a(n5739_1), .b(n5738) );
na02f01  g0253 ( .o(n5741), .a(n5740), .b(n5697) );
no02f01  g0254 ( .o(n5742), .a(n5740), .b(_net_9421) );
no02f01  g0255 ( .o(n5743), .a(n5742), .b(n5697) );
ao22f01  g0256 ( .o(n5744_1), .a(n5743), .b(x1743), .c(n5742), .d(_net_9414) );
oa12f01  g0257 ( .o(n528), .a(n5744_1), .b(n5741), .c(n5737) );
no02f01  g0258 ( .o(n5746), .a(_net_10118), .b(_net_10119) );
in01f01  g0259 ( .o(n5747), .a(n5746) );
ao12f01  g0260 ( .o(n5748_1), .a(_net_10116), .b(_net_10114), .c(_net_10115) );
in01f01  g0261 ( .o(n5749), .a(n5748_1) );
no02f01  g0262 ( .o(n5750), .a(n5749), .b(_net_10117) );
in01f01  g0263 ( .o(n5751), .a(n5750) );
no02f01  g0264 ( .o(n5752), .a(n5751), .b(n5747) );
in01f01  g0265 ( .o(n5753_1), .a(n5752) );
no02f01  g0266 ( .o(n5754), .a(n5753_1), .b(_net_10120) );
in01f01  g0267 ( .o(n5755), .a(n5754) );
no02f01  g0268 ( .o(n5756), .a(n5755), .b(_net_10121) );
in01f01  g0269 ( .o(n5757), .a(n5756) );
no02f01  g0270 ( .o(n5758_1), .a(n5757), .b(_net_10122) );
in01f01  g0271 ( .o(n5759), .a(n5758_1) );
no02f01  g0272 ( .o(n5760), .a(n5759), .b(_net_10123) );
in01f01  g0273 ( .o(n5761), .a(n5760) );
no02f01  g0274 ( .o(n5762), .a(n5761), .b(_net_10124) );
in01f01  g0275 ( .o(n5763_1), .a(n5762) );
na02f01  g0276 ( .o(n5764), .a(n5761), .b(_net_10124) );
na02f01  g0277 ( .o(n533), .a(n5764), .b(n5763_1) );
in01f01  g0278 ( .o(n5766), .a(_net_10312) );
no02f01  g0279 ( .o(n5767), .a(n5558), .b(x6577) );
no02f01  g0280 ( .o(n5768_1), .a(n5767), .b(n5658) );
no02f01  g0281 ( .o(n5769), .a(n5689), .b(n5658) );
no02f01  g0282 ( .o(n5770), .a(n5769), .b(n5768_1) );
in01f01  g0283 ( .o(n5771), .a(n5767) );
no02f01  g0284 ( .o(n5772), .a(n5771), .b(n5658) );
in01f01  g0285 ( .o(n5773_1), .a(n5772) );
no02f01  g0286 ( .o(n5774), .a(n5773_1), .b(n5690_1) );
ao12f01  g0287 ( .o(n5775), .a(n5658), .b(n5774), .c(x5647) );
oa12f01  g0288 ( .o(n538), .a(n5775), .b(n5770), .c(n5766) );
no02f01  g0289 ( .o(n5777_1), .a(net_194), .b(_net_9744) );
in01f01  g0290 ( .o(n5778), .a(_net_9744) );
in01f01  g0291 ( .o(n5779), .a(net_194) );
no02f01  g0292 ( .o(n5780), .a(n5779), .b(n5778) );
no02f01  g0293 ( .o(n5781), .a(_net_193), .b(_net_9743) );
in01f01  g0294 ( .o(n5782_1), .a(_net_9743) );
in01f01  g0295 ( .o(n5783), .a(_net_193) );
no02f01  g0296 ( .o(n5784), .a(n5783), .b(n5782_1) );
oa22f01  g0297 ( .o(n5785), .a(n5784), .b(n5781), .c(n5780), .d(n5777_1) );
in01f01  g0298 ( .o(n5786), .a(_net_9745) );
in01f01  g0299 ( .o(n5787_1), .a(net_195) );
no02f01  g0300 ( .o(n5788), .a(n5787_1), .b(n5786) );
no02f01  g0301 ( .o(n5789), .a(net_195), .b(_net_9745) );
no02f01  g0302 ( .o(n5790), .a(_net_9746), .b(net_196) );
in01f01  g0303 ( .o(n5791), .a(net_196) );
in01f01  g0304 ( .o(n5792_1), .a(_net_9746) );
no02f01  g0305 ( .o(n5793), .a(n5792_1), .b(n5791) );
oa22f01  g0306 ( .o(n5794), .a(n5793), .b(n5790), .c(n5789), .d(n5788) );
no02f01  g0307 ( .o(n3141), .a(n5794), .b(n5785) );
no02f01  g0308 ( .o(n5796), .a(_net_9845), .b(net_196) );
in01f01  g0309 ( .o(n5797_1), .a(_net_9845) );
no02f01  g0310 ( .o(n5798), .a(n5797_1), .b(n5791) );
in01f01  g0311 ( .o(n5799), .a(_net_9844) );
no02f01  g0312 ( .o(n5800), .a(n5787_1), .b(n5799) );
no02f01  g0313 ( .o(n5801), .a(net_195), .b(_net_9844) );
oa22f01  g0314 ( .o(n5802_1), .a(n5801), .b(n5800), .c(n5798), .d(n5796) );
in01f01  g0315 ( .o(n5803), .a(_net_9842) );
no02f01  g0316 ( .o(n5804), .a(n5803), .b(n5783) );
no02f01  g0317 ( .o(n5805), .a(_net_9842), .b(_net_193) );
in01f01  g0318 ( .o(n5806), .a(_net_9843) );
no02f01  g0319 ( .o(n5807_1), .a(n5806), .b(n5779) );
no02f01  g0320 ( .o(n5808), .a(_net_9843), .b(net_194) );
oa22f01  g0321 ( .o(n5809), .a(n5808), .b(n5807_1), .c(n5805), .d(n5804) );
no02f01  g0322 ( .o(n7557), .a(n5809), .b(n5802_1) );
no02f01  g0323 ( .o(n5811), .a(_net_9944), .b(net_196) );
in01f01  g0324 ( .o(n5812_1), .a(_net_9944) );
no02f01  g0325 ( .o(n5813), .a(n5812_1), .b(n5791) );
no02f01  g0326 ( .o(n5814), .a(net_195), .b(_net_9943) );
in01f01  g0327 ( .o(n5815_1), .a(_net_9943) );
no02f01  g0328 ( .o(n5816), .a(n5787_1), .b(n5815_1) );
oa22f01  g0329 ( .o(n5817), .a(n5816), .b(n5814), .c(n5813), .d(n5811) );
in01f01  g0330 ( .o(n5818), .a(_net_9941) );
no02f01  g0331 ( .o(n5819), .a(n5783), .b(n5818) );
no02f01  g0332 ( .o(n5820_1), .a(_net_193), .b(_net_9941) );
in01f01  g0333 ( .o(n5821), .a(_net_9942) );
no02f01  g0334 ( .o(n5822), .a(n5821), .b(n5779) );
no02f01  g0335 ( .o(n5823), .a(_net_9942), .b(net_194) );
oa22f01  g0336 ( .o(n5824), .a(n5823), .b(n5822), .c(n5820_1), .d(n5819) );
no02f01  g0337 ( .o(n7590), .a(n5824), .b(n5817) );
no02f01  g0338 ( .o(n5826), .a(_net_10043), .b(net_196) );
in01f01  g0339 ( .o(n5827), .a(_net_10043) );
no02f01  g0340 ( .o(n5828), .a(n5827), .b(n5791) );
in01f01  g0341 ( .o(n5829), .a(_net_10042) );
no02f01  g0342 ( .o(n5830_1), .a(n5787_1), .b(n5829) );
no02f01  g0343 ( .o(n5831), .a(net_195), .b(_net_10042) );
oa22f01  g0344 ( .o(n5832), .a(n5831), .b(n5830_1), .c(n5828), .d(n5826) );
in01f01  g0345 ( .o(n5833), .a(_net_10040) );
no02f01  g0346 ( .o(n5834), .a(n5783), .b(n5833) );
no02f01  g0347 ( .o(n5835_1), .a(_net_193), .b(_net_10040) );
in01f01  g0348 ( .o(n5836), .a(_net_10041) );
no02f01  g0349 ( .o(n5837), .a(n5836), .b(n5779) );
no02f01  g0350 ( .o(n5838), .a(_net_10041), .b(net_194) );
oa22f01  g0351 ( .o(n5839_1), .a(n5838), .b(n5837), .c(n5835_1), .d(n5834) );
no02f01  g0352 ( .o(n2794), .a(n5839_1), .b(n5832) );
no04f01  g0353 ( .o(n5841), .a(n2794), .b(n7590), .c(n7557), .d(n3141) );
no02f01  g0354 ( .o(n5842), .a(n5794), .b(n5785) );
ao22f01  g0355 ( .o(n5843), .a(n5842), .b(net_9678), .c(n5841), .d(net_116) );
no02f01  g0356 ( .o(n5844_1), .a(n7557), .b(n3141) );
in01f01  g0357 ( .o(n5845), .a(n7590) );
na03f01  g0358 ( .o(n5846), .a(n2794), .b(n5845), .c(n5844_1) );
no02f01  g0359 ( .o(n5847), .a(n5841), .b(n5846) );
na02f01  g0360 ( .o(n5848), .a(n5847), .b(net_9975) );
no03f01  g0361 ( .o(n5849_1), .a(n5845), .b(n7557), .c(n3141) );
no03f01  g0362 ( .o(n5850), .a(n5809), .b(n5802_1), .c(n3141) );
ao22f01  g0363 ( .o(n5851), .a(n5850), .b(net_9777), .c(n5849_1), .d(net_9876) );
na03f01  g0364 ( .o(n543), .a(n5851), .b(n5848), .c(n5843) );
in01f01  g0365 ( .o(n5853_1), .a(net_9513) );
no02f01  g0366 ( .o(n5854), .a(n5853_1), .b(_net_9250) );
in01f01  g0367 ( .o(n5855), .a(net_9539) );
no03f01  g0368 ( .o(n5856), .a(n5855), .b(_net_9515), .c(_net_9250) );
no02f01  g0369 ( .o(n5857), .a(n5856), .b(n5854) );
in01f01  g0370 ( .o(n5858_1), .a(net_9531) );
no02f01  g0371 ( .o(n5859), .a(n5858_1), .b(n5658) );
na03f01  g0372 ( .o(n5860), .a(n5859), .b(n5857), .c(net_9538) );
in01f01  g0373 ( .o(n5861), .a(net_9538) );
ao12f01  g0374 ( .o(n5862), .a(_net_9250), .b(n5489), .c(n5861) );
na03f01  g0375 ( .o(n5863_1), .a(n5862), .b(_net_9537), .c(x6599) );
in01f01  g0376 ( .o(n5864), .a(_net_9532) );
no02f01  g0377 ( .o(n5865), .a(n5864), .b(n5658) );
in01f01  g0378 ( .o(n5866), .a(n5865) );
na02f01  g0379 ( .o(n5867), .a(_net_9536), .b(x6599) );
na02f01  g0380 ( .o(n5868_1), .a(n5867), .b(n5866) );
na02f01  g0381 ( .o(n5869), .a(n5489), .b(net_9538) );
no02f01  g0382 ( .o(n5870), .a(n5869), .b(_net_9250) );
na02f01  g0383 ( .o(n5871), .a(net_9535), .b(x6599) );
no02f01  g0384 ( .o(n5872), .a(n5871), .b(n5869) );
ao12f01  g0385 ( .o(n5873_1), .a(n5872), .b(n5870), .c(n5868_1) );
no02f01  g0386 ( .o(n5874), .a(_net_9250), .b(n5861) );
no02f01  g0387 ( .o(n5875), .a(n5861), .b(n5658) );
in01f01  g0388 ( .o(n5876), .a(n5875) );
na03f01  g0389 ( .o(n5877), .a(_net_8869), .b(_net_9040), .c(_net_9383) );
no02f01  g0390 ( .o(n5878_1), .a(n5877), .b(n5739_1) );
no02f01  g0391 ( .o(n5879), .a(n5878_1), .b(n5876) );
no02f01  g0392 ( .o(n5880), .a(_net_9250), .b(_net_9530) );
in01f01  g0393 ( .o(n5881), .a(n5880) );
no02f01  g0394 ( .o(n5882), .a(n5881), .b(n5861) );
in01f01  g0395 ( .o(n5883_1), .a(net_9542) );
in01f01  g0396 ( .o(n5884), .a(net_9534) );
no02f01  g0397 ( .o(n5885), .a(n5884), .b(n5658) );
in01f01  g0398 ( .o(n5886), .a(n5885) );
no02f01  g0399 ( .o(n5887), .a(n5886), .b(net_9544) );
na02f01  g0400 ( .o(n5888_1), .a(n5887), .b(n5883_1) );
in01f01  g0401 ( .o(n5889), .a(net_9533) );
no02f01  g0402 ( .o(n5890), .a(n5889), .b(n5658) );
in01f01  g0403 ( .o(n5891), .a(n5890) );
oa12f01  g0404 ( .o(n5892), .a(n5888_1), .b(n5891), .c(_net_9503) );
ao22f01  g0405 ( .o(n5893_1), .a(n5892), .b(n5874), .c(n5882), .d(n5879) );
na04f01  g0406 ( .o(n548), .a(n5893_1), .b(n5873_1), .c(n5863_1), .d(n5860) );
in01f01  g0407 ( .o(n5895), .a(net_9940) );
oa22f01  g0408 ( .o(n553), .a(n5694), .b(n5895), .c(n5692), .d(n5591) );
in01f01  g0409 ( .o(n5897), .a(_net_10029) );
no02f01  g0410 ( .o(n5898_1), .a(n5549), .b(n5564) );
in01f01  g0411 ( .o(n5899), .a(n5898_1) );
no03f01  g0412 ( .o(n5900), .a(n5899), .b(n5666_1), .c(n5631) );
in01f01  g0413 ( .o(n5901), .a(n5900) );
no02f01  g0414 ( .o(n5902), .a(n5901), .b(n5664) );
in01f01  g0415 ( .o(n5903_1), .a(n5902) );
no02f01  g0416 ( .o(n5904), .a(n5903_1), .b(n5686) );
na02f01  g0417 ( .o(n5905), .a(n5904), .b(x6599) );
in01f01  g0418 ( .o(n5906), .a(n5904) );
na02f01  g0419 ( .o(n5907), .a(n5906), .b(x6599) );
oa22f01  g0420 ( .o(n563), .a(n5907), .b(n5897), .c(n5905), .d(n5561) );
in01f01  g0421 ( .o(n5909), .a(net_10299) );
in01f01  g0422 ( .o(n5910), .a(net_10293) );
na02f01  g0423 ( .o(n5911), .a(n5910), .b(x6599) );
na02f01  g0424 ( .o(n5912), .a(net_263), .b(net_10280) );
ao12f01  g0425 ( .o(n568), .a(n5911), .b(n5912), .c(n5909) );
in01f01  g0426 ( .o(n5914), .a(net_9273) );
no02f01  g0427 ( .o(n573), .a(_net_9268), .b(n5914) );
in01f01  g0428 ( .o(n5916), .a(_net_168) );
in01f01  g0429 ( .o(n5917_1), .a(_net_8828) );
in01f01  g0430 ( .o(n5918), .a(_net_188) );
ao12f01  g0431 ( .o(n5919), .a(_net_187), .b(n5918), .c(n5917_1) );
in01f01  g0432 ( .o(n5920), .a(_net_180) );
no02f01  g0433 ( .o(n5921_1), .a(_net_188), .b(_net_187) );
no02f01  g0434 ( .o(n5922), .a(n5921_1), .b(n5920) );
na02f01  g0435 ( .o(n5923), .a(n5922), .b(n5919) );
in01f01  g0436 ( .o(n5924), .a(n5923) );
oa12f01  g0437 ( .o(n5925), .a(n5918), .b(_net_9572), .c(_net_187) );
in01f01  g0438 ( .o(n5926_1), .a(n5925) );
na02f01  g0439 ( .o(n5927), .a(n5926_1), .b(n5923) );
in01f01  g0440 ( .o(n5928), .a(n5927) );
in01f01  g0441 ( .o(n5929), .a(n5922) );
in01f01  g0442 ( .o(n5930), .a(_net_9572) );
in01f01  g0443 ( .o(n5931_1), .a(n5921_1) );
no02f01  g0444 ( .o(n5932), .a(n5931_1), .b(n5930) );
no02f01  g0445 ( .o(n5933), .a(_net_9562), .b(_net_191) );
no03f01  g0446 ( .o(n5934), .a(n5933), .b(n5921_1), .c(_net_9565) );
oa12f01  g0447 ( .o(n5935_1), .a(n5929), .b(n5934), .c(n5932) );
in01f01  g0448 ( .o(n5936), .a(_net_153) );
no02f01  g0449 ( .o(n5937), .a(n5935_1), .b(n5936) );
ao12f01  g0450 ( .o(n5938), .a(n5937), .b(n5935_1), .c(_net_119) );
in01f01  g0451 ( .o(n5939_1), .a(_net_154) );
no02f01  g0452 ( .o(n5940), .a(n5935_1), .b(n5939_1) );
ao12f01  g0453 ( .o(n5941), .a(n5940), .b(n5935_1), .c(_net_120) );
ao22f01  g0454 ( .o(n5942), .a(n5941), .b(_net_170), .c(n5938), .d(_net_169) );
in01f01  g0455 ( .o(n5943), .a(_net_152) );
no02f01  g0456 ( .o(n5944_1), .a(n5935_1), .b(n5943) );
ao12f01  g0457 ( .o(n5945), .a(n5944_1), .b(n5935_1), .c(_net_118) );
in01f01  g0458 ( .o(n5946), .a(_net_151) );
no02f01  g0459 ( .o(n5947), .a(n5935_1), .b(n5946) );
ao12f01  g0460 ( .o(n5948), .a(n5947), .b(n5935_1), .c(_net_117) );
ao22f01  g0461 ( .o(n5949_1), .a(n5948), .b(_net_167), .c(n5945), .d(_net_168) );
no02f01  g0462 ( .o(n5950), .a(n5945), .b(_net_168) );
oa12f01  g0463 ( .o(n5951), .a(n5942), .b(n5950), .c(n5949_1) );
no03f01  g0464 ( .o(n5952), .a(n5941), .b(n5938), .c(_net_169) );
no03f01  g0465 ( .o(n5953), .a(n5938), .b(_net_169), .c(_net_170) );
no02f01  g0466 ( .o(n5954_1), .a(n5941), .b(_net_170) );
no03f01  g0467 ( .o(n5955), .a(n5954_1), .b(n5953), .c(n5952) );
in01f01  g0468 ( .o(n5956), .a(_net_158) );
no02f01  g0469 ( .o(n5957), .a(n5935_1), .b(n5956) );
ao12f01  g0470 ( .o(n5958), .a(n5957), .b(n5935_1), .c(_net_124) );
in01f01  g0471 ( .o(n5959_1), .a(_net_157) );
no02f01  g0472 ( .o(n5960), .a(n5935_1), .b(n5959_1) );
ao12f01  g0473 ( .o(n5961), .a(n5960), .b(n5935_1), .c(_net_123) );
ao22f01  g0474 ( .o(n5962), .a(n5961), .b(_net_173), .c(n5958), .d(_net_174) );
in01f01  g0475 ( .o(n5963), .a(_net_155) );
no02f01  g0476 ( .o(n5964_1), .a(n5935_1), .b(n5963) );
ao12f01  g0477 ( .o(n5965), .a(n5964_1), .b(n5935_1), .c(_net_121) );
in01f01  g0478 ( .o(n5966), .a(_net_156) );
no02f01  g0479 ( .o(n5967), .a(n5935_1), .b(n5966) );
ao12f01  g0480 ( .o(n5968), .a(n5967), .b(n5935_1), .c(_net_122) );
ao22f01  g0481 ( .o(n5969_1), .a(n5968), .b(_net_172), .c(n5965), .d(_net_171) );
na02f01  g0482 ( .o(n5970), .a(n5969_1), .b(n5962) );
ao12f01  g0483 ( .o(n5971), .a(n5970), .b(n5955), .c(n5951) );
no03f01  g0484 ( .o(n5972), .a(n5968), .b(n5965), .c(_net_171) );
no03f01  g0485 ( .o(n5973), .a(n5965), .b(_net_171), .c(_net_172) );
oa12f01  g0486 ( .o(n5974_1), .a(n5962), .b(n5973), .c(n5972) );
in01f01  g0487 ( .o(n5975), .a(_net_172) );
in01f01  g0488 ( .o(n5976), .a(n5968) );
na03f01  g0489 ( .o(n5977), .a(n5976), .b(n5962), .c(n5975) );
no03f01  g0490 ( .o(n5978_1), .a(n5961), .b(_net_173), .c(_net_174) );
no03f01  g0491 ( .o(n5979), .a(n5961), .b(n5958), .c(_net_173) );
no02f01  g0492 ( .o(n5980), .a(n5958), .b(_net_174) );
no03f01  g0493 ( .o(n5981), .a(n5980), .b(n5979), .c(n5978_1) );
na03f01  g0494 ( .o(n5982), .a(n5981), .b(n5977), .c(n5974_1) );
in01f01  g0495 ( .o(n5983_1), .a(_net_177) );
in01f01  g0496 ( .o(n5984), .a(_net_161) );
no02f01  g0497 ( .o(n5985), .a(n5935_1), .b(n5984) );
ao12f01  g0498 ( .o(n5986), .a(n5985), .b(n5935_1), .c(_net_127) );
in01f01  g0499 ( .o(n5987), .a(n5986) );
no02f01  g0500 ( .o(n5988_1), .a(n5987), .b(n5983_1) );
in01f01  g0501 ( .o(n5989), .a(_net_175) );
in01f01  g0502 ( .o(n5990), .a(_net_176) );
in01f01  g0503 ( .o(n5991), .a(_net_160) );
no02f01  g0504 ( .o(n5992), .a(n5935_1), .b(n5991) );
ao12f01  g0505 ( .o(n5993_1), .a(n5992), .b(n5935_1), .c(_net_126) );
in01f01  g0506 ( .o(n5994), .a(n5993_1) );
in01f01  g0507 ( .o(n5995), .a(_net_159) );
no02f01  g0508 ( .o(n5996), .a(n5935_1), .b(n5995) );
ao12f01  g0509 ( .o(n5997), .a(n5996), .b(n5935_1), .c(_net_125) );
in01f01  g0510 ( .o(n5998_1), .a(n5997) );
oa22f01  g0511 ( .o(n5999), .a(n5998_1), .b(n5989), .c(n5994), .d(n5990) );
no02f01  g0512 ( .o(n6000), .a(n5999), .b(n5988_1) );
oa12f01  g0513 ( .o(n6001_1), .a(n6000), .b(n5982), .c(n5971) );
in01f01  g0514 ( .o(n6002), .a(n6001_1) );
no03f01  g0515 ( .o(n6003), .a(n5997), .b(_net_176), .c(_net_175) );
no03f01  g0516 ( .o(n6004), .a(n5997), .b(n5993_1), .c(_net_175) );
no02f01  g0517 ( .o(n6005_1), .a(n5993_1), .b(_net_176) );
no02f01  g0518 ( .o(n6006), .a(n5986), .b(_net_177) );
no04f01  g0519 ( .o(n6007), .a(n6006), .b(n6005_1), .c(n6004), .d(n6003) );
na02f01  g0520 ( .o(n6008), .a(n5935_1), .b(_net_128) );
in01f01  g0521 ( .o(n6009_1), .a(n5935_1) );
na02f01  g0522 ( .o(n6010), .a(n6009_1), .b(_net_162) );
na02f01  g0523 ( .o(n6011), .a(n6010), .b(n6008) );
na02f01  g0524 ( .o(n6012), .a(n5935_1), .b(_net_130) );
na02f01  g0525 ( .o(n6013_1), .a(n6009_1), .b(_net_164) );
na02f01  g0526 ( .o(n6014), .a(n6013_1), .b(n6012) );
na02f01  g0527 ( .o(n6015), .a(n5935_1), .b(_net_129) );
na02f01  g0528 ( .o(n6016), .a(n6009_1), .b(_net_163) );
na02f01  g0529 ( .o(n6017), .a(n6016), .b(n6015) );
no03f01  g0530 ( .o(n6018_1), .a(n6017), .b(n6014), .c(n6011) );
oa12f01  g0531 ( .o(n6019), .a(n6018_1), .b(n6007), .c(n5988_1) );
no02f01  g0532 ( .o(n6020), .a(n6019), .b(n6002) );
in01f01  g0533 ( .o(n6021), .a(n6020) );
ao12f01  g0534 ( .o(n6022), .a(n5924), .b(n6021), .c(n5928) );
na02f01  g0535 ( .o(n6023_1), .a(n5935_1), .b(_net_118) );
oa12f01  g0536 ( .o(n6024), .a(n6023_1), .b(n5935_1), .c(n5943) );
in01f01  g0537 ( .o(n6025), .a(_net_9291) );
na02f01  g0538 ( .o(n6026), .a(n5925), .b(n5923) );
no02f01  g0539 ( .o(n6027), .a(n6026), .b(n6025) );
no02f01  g0540 ( .o(n6028_1), .a(n6021), .b(n5927) );
ao12f01  g0541 ( .o(n6029), .a(n6027), .b(n6028_1), .c(n6024) );
oa12f01  g0542 ( .o(n578), .a(n6029), .b(n6022), .c(n5916) );
in01f01  g0543 ( .o(n6031), .a(_net_132) );
in01f01  g0544 ( .o(n6032), .a(n5770) );
na04f01  g0545 ( .o(n6033_1), .a(n6032), .b(_net_133), .c(net_10385), .d(n6031) );
na03f01  g0546 ( .o(n6034), .a(n6032), .b(net_10385), .c(_net_132) );
no02f01  g0547 ( .o(n6035), .a(n5774), .b(n5658) );
na03f01  g0548 ( .o(n6036), .a(n6035), .b(n6034), .c(n6033_1) );
in01f01  g0549 ( .o(n6037_1), .a(n6036) );
no02f01  g0550 ( .o(n6038), .a(n6037_1), .b(n6033_1) );
na02f01  g0551 ( .o(n6039), .a(n6038), .b(net_240) );
na02f01  g0552 ( .o(n6040), .a(n6036), .b(n5658) );
na02f01  g0553 ( .o(n6041), .a(n6037_1), .b(net_9869) );
no02f01  g0554 ( .o(n6042_1), .a(n6037_1), .b(n6034) );
in01f01  g0555 ( .o(n6043), .a(n5774) );
no02f01  g0556 ( .o(n6044), .a(n6037_1), .b(n6043) );
ao22f01  g0557 ( .o(n6045), .a(n6044), .b(x5548), .c(n6042_1), .d(_net_10314) );
na04f01  g0558 ( .o(n583), .a(n6045), .b(n6041), .c(n6040), .d(n6039) );
no02f01  g0559 ( .o(n6047_1), .a(n5902), .b(n5658) );
no02f01  g0560 ( .o(n6048), .a(n6047_1), .b(n5768_1) );
in01f01  g0561 ( .o(n6049), .a(n6048) );
na04f01  g0562 ( .o(n6050), .a(n6049), .b(_net_133), .c(n6031), .d(net_10490) );
na03f01  g0563 ( .o(n6051), .a(n6049), .b(_net_132), .c(net_10490) );
no02f01  g0564 ( .o(n6052_1), .a(n5903_1), .b(n5773_1) );
no02f01  g0565 ( .o(n6053), .a(n6052_1), .b(n5658) );
na03f01  g0566 ( .o(n6054), .a(n6053), .b(n6051), .c(n6050) );
in01f01  g0567 ( .o(n6055), .a(n6054) );
no02f01  g0568 ( .o(n6056), .a(n6055), .b(n6050) );
na02f01  g0569 ( .o(n6057_1), .a(n6056), .b(net_262) );
na02f01  g0570 ( .o(n6058), .a(n6054), .b(n5658) );
na02f01  g0571 ( .o(n6059), .a(n6055), .b(net_9990) );
no02f01  g0572 ( .o(n6060), .a(n6055), .b(n6051) );
in01f01  g0573 ( .o(n6061), .a(n6052_1) );
no02f01  g0574 ( .o(n6062_1), .a(n6055), .b(n6061) );
ao22f01  g0575 ( .o(n6063), .a(n6062_1), .b(x3889), .c(n6060), .d(_net_10441) );
na04f01  g0576 ( .o(n588), .a(n6063), .b(n6059), .c(n6058), .d(n6057_1) );
na02f01  g0577 ( .o(n6065), .a(n5877), .b(n5738) );
in01f01  g0578 ( .o(n6066), .a(n6065) );
in01f01  g0579 ( .o(n6067_1), .a(_net_8955) );
no02f01  g0580 ( .o(n6068), .a(n6067_1), .b(_net_9062) );
no02f01  g0581 ( .o(n6069), .a(n6068), .b(n5699) );
na03f01  g0582 ( .o(n6070), .a(n5877), .b(_net_8955), .c(n5738) );
oa12f01  g0583 ( .o(n6071), .a(n6070), .b(n6069), .c(n6066) );
na03f01  g0584 ( .o(n6072_1), .a(n5877), .b(_net_9062), .c(n5738) );
in01f01  g0585 ( .o(n6073), .a(n6072_1) );
ao12f01  g0586 ( .o(n6074), .a(_net_9062), .b(n5877), .c(n5738) );
no02f01  g0587 ( .o(n6075), .a(n6074), .b(n6073) );
in01f01  g0588 ( .o(n6076), .a(_net_9388) );
ao12f01  g0589 ( .o(n6077_1), .a(n6076), .b(_net_8955), .c(_net_9062) );
no02f01  g0590 ( .o(n6078), .a(n5739_1), .b(_net_9388) );
no02f01  g0591 ( .o(n6079), .a(n6078), .b(n6077_1) );
na03f01  g0592 ( .o(n6080), .a(n5877), .b(_net_9388), .c(n5738) );
oa12f01  g0593 ( .o(n6081), .a(n6080), .b(n6079), .c(n6066) );
na04f01  g0594 ( .o(n6082_1), .a(n6081), .b(n6075), .c(n6071), .d(net_9486) );
in01f01  g0595 ( .o(n6083), .a(n6074) );
na02f01  g0596 ( .o(n6084), .a(n6083), .b(n6072_1) );
na04f01  g0597 ( .o(n6085), .a(n6081), .b(n6084), .c(n6071), .d(net_9494) );
na02f01  g0598 ( .o(n6086), .a(n6067_1), .b(_net_9062) );
na02f01  g0599 ( .o(n6087_1), .a(_net_8955), .b(n5698) );
ao22f01  g0600 ( .o(n6088), .a(n6087_1), .b(n6086), .c(n5877), .d(n5738) );
ao12f01  g0601 ( .o(n6089), .a(n6088), .b(n6066), .c(_net_8955) );
na04f01  g0602 ( .o(n6090), .a(n6081), .b(n6075), .c(n6089), .d(net_9470) );
na04f01  g0603 ( .o(n6091_1), .a(n6081), .b(n6084), .c(n6089), .d(net_9478) );
na04f01  g0604 ( .o(n6092), .a(n6091_1), .b(n6090), .c(n6085), .d(n6082_1) );
na02f01  g0605 ( .o(n6093), .a(n5739_1), .b(_net_9388) );
na03f01  g0606 ( .o(n6094), .a(n6076), .b(_net_8955), .c(_net_9062) );
na02f01  g0607 ( .o(n6095_1), .a(n6094), .b(n6093) );
in01f01  g0608 ( .o(n6096), .a(n6080) );
ao12f01  g0609 ( .o(n6097), .a(n6096), .b(n6095_1), .c(n6065) );
na04f01  g0610 ( .o(n6098), .a(n6097), .b(n6075), .c(n6071), .d(net_9454) );
na04f01  g0611 ( .o(n6099_1), .a(n6097), .b(n6084), .c(n6071), .d(net_9462) );
na04f01  g0612 ( .o(n6100), .a(n6097), .b(n6075), .c(n6089), .d(net_9438) );
na04f01  g0613 ( .o(n6101), .a(n6097), .b(n6084), .c(n6089), .d(net_9446) );
na04f01  g0614 ( .o(n6102_1), .a(n6101), .b(n6100), .c(n6099_1), .d(n6098) );
no02f01  g0615 ( .o(n6103), .a(n6102_1), .b(n6092) );
in01f01  g0616 ( .o(n6104), .a(_net_9363) );
no02f01  g0617 ( .o(n6105), .a(n6104), .b(_net_9377) );
in01f01  g0618 ( .o(n6106), .a(_net_9377) );
no02f01  g0619 ( .o(n6107_1), .a(_net_9363), .b(n6106) );
no02f01  g0620 ( .o(n6108), .a(n6107_1), .b(n6105) );
no02f01  g0621 ( .o(n6109), .a(n6108), .b(n6103) );
in01f01  g0622 ( .o(n6110), .a(net_9486) );
no04f01  g0623 ( .o(n6111_1), .a(n6097), .b(n6084), .c(n6089), .d(n6110) );
in01f01  g0624 ( .o(n6112), .a(net_9494) );
no04f01  g0625 ( .o(n6113), .a(n6097), .b(n6075), .c(n6089), .d(n6112) );
in01f01  g0626 ( .o(n6114), .a(net_9470) );
no04f01  g0627 ( .o(n6115), .a(n6097), .b(n6084), .c(n6071), .d(n6114) );
in01f01  g0628 ( .o(n6116_1), .a(net_9478) );
no04f01  g0629 ( .o(n6117), .a(n6097), .b(n6075), .c(n6071), .d(n6116_1) );
no04f01  g0630 ( .o(n6118), .a(n6117), .b(n6115), .c(n6113), .d(n6111_1) );
in01f01  g0631 ( .o(n6119), .a(net_9454) );
no04f01  g0632 ( .o(n6120), .a(n6081), .b(n6084), .c(n6089), .d(n6119) );
in01f01  g0633 ( .o(n6121_1), .a(net_9462) );
no04f01  g0634 ( .o(n6122), .a(n6081), .b(n6075), .c(n6089), .d(n6121_1) );
in01f01  g0635 ( .o(n6123), .a(net_9438) );
no04f01  g0636 ( .o(n6124), .a(n6081), .b(n6084), .c(n6071), .d(n6123) );
in01f01  g0637 ( .o(n6125), .a(net_9446) );
no04f01  g0638 ( .o(n6126_1), .a(n6081), .b(n6075), .c(n6071), .d(n6125) );
no04f01  g0639 ( .o(n6127), .a(n6126_1), .b(n6124), .c(n6122), .d(n6120) );
na02f01  g0640 ( .o(n6128), .a(n6127), .b(n6118) );
in01f01  g0641 ( .o(n6129), .a(n6108) );
no02f01  g0642 ( .o(n6130), .a(_net_9514), .b(_net_9515) );
no02f01  g0643 ( .o(n6131_1), .a(n6130), .b(_net_9378) );
in01f01  g0644 ( .o(n6132), .a(n5877) );
in01f01  g0645 ( .o(n6133), .a(_net_9378) );
no03f01  g0646 ( .o(n6134), .a(net_9379), .b(n6133), .c(_net_8825) );
in01f01  g0647 ( .o(n6135), .a(_net_9383) );
in01f01  g0648 ( .o(n6136_1), .a(_net_9040) );
in01f01  g0649 ( .o(n6137), .a(_net_8869) );
in01f01  g0650 ( .o(n7446), .a(n6130) );
no03f01  g0651 ( .o(n6139), .a(n7446), .b(n6137), .c(n6136_1) );
in01f01  g0652 ( .o(n6140), .a(n6139) );
no02f01  g0653 ( .o(n6141_1), .a(n6140), .b(n6135) );
in01f01  g0654 ( .o(n6142), .a(_net_9384) );
no02f01  g0655 ( .o(n6143), .a(n6142), .b(_net_9040) );
no02f01  g0656 ( .o(n6144), .a(n6143), .b(_net_9386) );
in01f01  g0657 ( .o(n6145_1), .a(n6144) );
no02f01  g0658 ( .o(n6146), .a(n6145_1), .b(n6141_1) );
ao12f01  g0659 ( .o(n6147), .a(n6134), .b(n6146), .c(n6132) );
no02f01  g0660 ( .o(n6148), .a(n6147), .b(n6131_1) );
oa12f01  g0661 ( .o(n6149), .a(n6148), .b(n6129), .c(n6128) );
ao12f01  g0662 ( .o(n6150_1), .a(n6131_1), .b(n6147), .c(_net_9371) );
oa12f01  g0663 ( .o(n593), .a(n6150_1), .b(n6149), .c(n6109) );
in01f01  g0664 ( .o(n6152), .a(net_10065) );
in01f01  g0665 ( .o(n6153), .a(_net_10090) );
in01f01  g0666 ( .o(n6154), .a(net_10058) );
na02f01  g0667 ( .o(n6155_1), .a(n6154), .b(x6599) );
ao12f01  g0668 ( .o(n598), .a(n6155_1), .b(n6153), .c(n6152) );
in01f01  g0669 ( .o(n6157), .a(_net_10104) );
no02f01  g0670 ( .o(n6158), .a(n5671_1), .b(n5658) );
no02f01  g0671 ( .o(n6159), .a(n6158), .b(n5768_1) );
no02f01  g0672 ( .o(n6160_1), .a(n5773_1), .b(n5672) );
ao12f01  g0673 ( .o(n6161), .a(n5658), .b(n6160_1), .c(x5548) );
oa12f01  g0674 ( .o(n603), .a(n6161), .b(n6159), .c(n6157) );
in01f01  g0675 ( .o(n6163), .a(_net_9839) );
no02f01  g0676 ( .o(n6164_1), .a(_net_133), .b(_net_132) );
in01f01  g0677 ( .o(n6165), .a(n6164_1) );
oa12f01  g0678 ( .o(n6166), .a(net_10280), .b(n6165), .c(_net_8829) );
in01f01  g0679 ( .o(n6167), .a(n6166) );
no03f01  g0680 ( .o(n6168), .a(n6167), .b(net_10304), .c(n6163) );
na02f01  g0681 ( .o(n6169_1), .a(n6168), .b(_net_10258) );
no02f01  g0682 ( .o(n6170), .a(_net_10257), .b(_net_10258) );
in01f01  g0683 ( .o(n6171), .a(_net_10258) );
in01f01  g0684 ( .o(n6172), .a(_net_10257) );
no02f01  g0685 ( .o(n6173_1), .a(n6172), .b(n6171) );
in01f01  g0686 ( .o(n6174), .a(net_10304) );
no02f01  g0687 ( .o(n6175), .a(n6174), .b(n6163) );
oa12f01  g0688 ( .o(n6176), .a(n6175), .b(n6173_1), .c(n6170) );
no03f01  g0689 ( .o(n6177_1), .a(n6166), .b(net_10304), .c(n6163) );
in01f01  g0690 ( .o(n6178), .a(_net_9828) );
no02f01  g0691 ( .o(n6179), .a(n6178), .b(n6171) );
in01f01  g0692 ( .o(n6180), .a(n6179) );
no02f01  g0693 ( .o(n6181_1), .a(_net_9828), .b(_net_10258) );
in01f01  g0694 ( .o(n6182), .a(n6181_1) );
in01f01  g0695 ( .o(n6183), .a(_net_9827) );
no02f01  g0696 ( .o(n6184), .a(n6172), .b(n6183) );
na03f01  g0697 ( .o(n6185), .a(n6184), .b(n6182), .c(n6180) );
in01f01  g0698 ( .o(n6186_1), .a(n6184) );
oa12f01  g0699 ( .o(n6187), .a(n6186_1), .b(n6181_1), .c(n6179) );
na03f01  g0700 ( .o(n6188), .a(n6187), .b(n6185), .c(n6177_1) );
na03f01  g0701 ( .o(n608), .a(n6188), .b(n6176), .c(n6169_1) );
no02f01  g0702 ( .o(n6190), .a(_net_9421), .b(n5489) );
in01f01  g0703 ( .o(n6191_1), .a(_net_269) );
in01f01  g0704 ( .o(n6192), .a(_net_267) );
na02f01  g0705 ( .o(n6193), .a(_net_266), .b(_net_265) );
no02f01  g0706 ( .o(n6194), .a(n6193), .b(n6192) );
na02f01  g0707 ( .o(n6195), .a(n6194), .b(_net_268) );
no02f01  g0708 ( .o(n6196_1), .a(n6195), .b(n6191_1) );
na02f01  g0709 ( .o(n6197), .a(n6196_1), .b(_net_270) );
no02f01  g0710 ( .o(n6198), .a(n6197), .b(n5528_1) );
na02f01  g0711 ( .o(n6199), .a(n6198), .b(_net_272) );
no04f01  g0712 ( .o(n6200), .a(n5643), .b(n5579), .c(n5522), .d(n5534) );
in01f01  g0713 ( .o(n6201_1), .a(n6200) );
no02f01  g0714 ( .o(n6202), .a(n6201_1), .b(n6199) );
in01f01  g0715 ( .o(n6203), .a(n6202) );
no02f01  g0716 ( .o(n6204), .a(n6203), .b(_net_277) );
no02f01  g0717 ( .o(n6205), .a(n6202), .b(n5509) );
oa12f01  g0718 ( .o(n6206_1), .a(n6190), .b(n6205), .c(n6204) );
in01f01  g0719 ( .o(n6207), .a(n6190) );
na02f01  g0720 ( .o(n6208), .a(n6207), .b(_net_277) );
na02f01  g0721 ( .o(n6209), .a(n6208), .b(n6206_1) );
na02f01  g0722 ( .o(n6210), .a(n6209), .b(_net_9434) );
in01f01  g0723 ( .o(n6211_1), .a(_net_9434) );
na03f01  g0724 ( .o(n6212), .a(n6208), .b(n6206_1), .c(n6211_1) );
na02f01  g0725 ( .o(n6213), .a(n6212), .b(n6210) );
in01f01  g0726 ( .o(n6214), .a(net_9435) );
na02f01  g0727 ( .o(n6215), .a(n6202), .b(_net_277) );
no02f01  g0728 ( .o(n6216_1), .a(n6215), .b(_net_278) );
in01f01  g0729 ( .o(n6217), .a(n6215) );
no02f01  g0730 ( .o(n6218), .a(n6217), .b(n5543) );
oa12f01  g0731 ( .o(n6219), .a(n6190), .b(n6218), .c(n6216_1) );
na02f01  g0732 ( .o(n6220), .a(n6207), .b(_net_278) );
na02f01  g0733 ( .o(n6221_1), .a(n6220), .b(n6219) );
na02f01  g0734 ( .o(n6222), .a(n6221_1), .b(n6214) );
na03f01  g0735 ( .o(n6223), .a(n6220), .b(n6219), .c(net_9435) );
na03f01  g0736 ( .o(n6224), .a(n6223), .b(n6222), .c(n6213) );
na02f01  g0737 ( .o(n6225), .a(n6198), .b(n5588) );
in01f01  g0738 ( .o(n6226_1), .a(n6225) );
no02f01  g0739 ( .o(n6227), .a(n6198), .b(n5588) );
oa12f01  g0740 ( .o(n6228), .a(n6190), .b(n6227), .c(n6226_1) );
na02f01  g0741 ( .o(n6229), .a(n6207), .b(_net_272) );
na02f01  g0742 ( .o(n6230), .a(n6229), .b(n6228) );
na02f01  g0743 ( .o(n6231_1), .a(n6230), .b(_net_9429) );
in01f01  g0744 ( .o(n6232), .a(_net_9429) );
na03f01  g0745 ( .o(n6233), .a(n6229), .b(n6228), .c(n6232) );
in01f01  g0746 ( .o(n6234), .a(_net_9428) );
no02f01  g0747 ( .o(n6235_1), .a(n6197), .b(_net_271) );
ao12f01  g0748 ( .o(n6236), .a(n5528_1), .b(n6196_1), .c(_net_270) );
oa12f01  g0749 ( .o(n6237), .a(n6190), .b(n6236), .c(n6235_1) );
oa12f01  g0750 ( .o(n6238), .a(n6237), .b(n6190), .c(n5528_1) );
in01f01  g0751 ( .o(n6239), .a(n6238) );
no02f01  g0752 ( .o(n6240_1), .a(n6239), .b(n6234) );
no02f01  g0753 ( .o(n6241), .a(n6238), .b(_net_9428) );
no03f01  g0754 ( .o(n6242), .a(n6195), .b(_net_270), .c(n6191_1) );
no02f01  g0755 ( .o(n6243), .a(n6196_1), .b(n5652) );
oa12f01  g0756 ( .o(n6244_1), .a(n6190), .b(n6243), .c(n6242) );
oa12f01  g0757 ( .o(n6245), .a(n6244_1), .b(n6190), .c(n5652) );
na02f01  g0758 ( .o(n6246), .a(n6245), .b(_net_9427) );
in01f01  g0759 ( .o(n6247), .a(_net_9427) );
in01f01  g0760 ( .o(n6248), .a(n6245) );
na02f01  g0761 ( .o(n6249_1), .a(n6248), .b(n6247) );
in01f01  g0762 ( .o(n6250), .a(_net_9424) );
no02f01  g0763 ( .o(n6251), .a(n6193), .b(_net_267) );
ao12f01  g0764 ( .o(n6252), .a(n6192), .b(_net_266), .c(_net_265) );
oa12f01  g0765 ( .o(n6253), .a(n6190), .b(n6252), .c(n6251) );
oa12f01  g0766 ( .o(n6254_1), .a(n6253), .b(n6190), .c(n6192) );
in01f01  g0767 ( .o(n6255), .a(n6254_1) );
no02f01  g0768 ( .o(n6256), .a(n6255), .b(n6250) );
no02f01  g0769 ( .o(n6257), .a(n6254_1), .b(_net_9424) );
no02f01  g0770 ( .o(n6258_1), .a(n6257), .b(n6256) );
in01f01  g0771 ( .o(n6259), .a(_net_9423) );
in01f01  g0772 ( .o(n6260), .a(_net_266) );
in01f01  g0773 ( .o(n6261), .a(_net_265) );
no02f01  g0774 ( .o(n6262), .a(_net_266), .b(n6261) );
no02f01  g0775 ( .o(n6263_1), .a(n6260), .b(_net_265) );
oa12f01  g0776 ( .o(n6264), .a(n6190), .b(n6263_1), .c(n6262) );
oa12f01  g0777 ( .o(n6265), .a(n6264), .b(n6190), .c(n6260) );
in01f01  g0778 ( .o(n6266), .a(n6265) );
no02f01  g0779 ( .o(n6267), .a(n6266), .b(n6259) );
no02f01  g0780 ( .o(n6268_1), .a(n6265), .b(_net_9423) );
no02f01  g0781 ( .o(n6269), .a(n6268_1), .b(n6267) );
no02f01  g0782 ( .o(n6270), .a(n6207), .b(_net_265) );
no02f01  g0783 ( .o(n6271), .a(n6190), .b(n6261) );
no02f01  g0784 ( .o(n6272_1), .a(n6271), .b(n6270) );
ao12f01  g0785 ( .o(n6273), .a(n5929), .b(n6272_1), .c(_net_9422) );
oa12f01  g0786 ( .o(n6274), .a(n6273), .b(n6272_1), .c(_net_9422) );
in01f01  g0787 ( .o(n6275), .a(net_9425) );
in01f01  g0788 ( .o(n6276), .a(_net_268) );
no03f01  g0789 ( .o(n6277_1), .a(n6193), .b(n6192), .c(_net_268) );
no02f01  g0790 ( .o(n6278), .a(n6194), .b(n6276) );
oa12f01  g0791 ( .o(n6279), .a(n6190), .b(n6278), .c(n6277_1) );
oa12f01  g0792 ( .o(n6280), .a(n6279), .b(n6190), .c(n6276) );
na02f01  g0793 ( .o(n6281), .a(n6280), .b(n6275) );
in01f01  g0794 ( .o(n6282_1), .a(n6280) );
na02f01  g0795 ( .o(n6283), .a(n6282_1), .b(net_9425) );
na02f01  g0796 ( .o(n6284), .a(n6283), .b(n6281) );
no04f01  g0797 ( .o(n6285), .a(n6284), .b(n6274), .c(n6269), .d(n6258_1) );
in01f01  g0798 ( .o(n6286), .a(net_9426) );
no02f01  g0799 ( .o(n6287_1), .a(n6195), .b(_net_269) );
ao12f01  g0800 ( .o(n6288), .a(n6191_1), .b(n6194), .c(_net_268) );
oa12f01  g0801 ( .o(n6289), .a(n6190), .b(n6288), .c(n6287_1) );
oa12f01  g0802 ( .o(n6290), .a(n6289), .b(n6190), .c(n6191_1) );
na02f01  g0803 ( .o(n6291), .a(n6290), .b(n6286) );
in01f01  g0804 ( .o(n6292_1), .a(n6290) );
na02f01  g0805 ( .o(n6293), .a(n6292_1), .b(net_9426) );
na03f01  g0806 ( .o(n6294), .a(n6293), .b(n6291), .c(n6285) );
ao12f01  g0807 ( .o(n6295), .a(n6294), .b(n6249_1), .c(n6246) );
oa12f01  g0808 ( .o(n6296), .a(n6295), .b(n6241), .c(n6240_1) );
ao12f01  g0809 ( .o(n6297_1), .a(n6296), .b(n6233), .c(n6231_1) );
no02f01  g0810 ( .o(n6298), .a(n6199), .b(_net_273) );
na02f01  g0811 ( .o(n6299), .a(n6199), .b(_net_273) );
in01f01  g0812 ( .o(n6300), .a(n6299) );
oa12f01  g0813 ( .o(n6301), .a(n6190), .b(n6300), .c(n6298) );
na02f01  g0814 ( .o(n6302_1), .a(n6207), .b(_net_273) );
ao12f01  g0815 ( .o(n6303), .a(net_9430), .b(n6302_1), .c(n6301) );
in01f01  g0816 ( .o(n6304), .a(net_9430) );
na02f01  g0817 ( .o(n6305), .a(n6302_1), .b(n6301) );
no02f01  g0818 ( .o(n6306_1), .a(n6305), .b(n6304) );
no02f01  g0819 ( .o(n6307), .a(n6306_1), .b(n6303) );
in01f01  g0820 ( .o(n6308), .a(net_9431) );
no02f01  g0821 ( .o(n6309), .a(n6199), .b(n5643) );
in01f01  g0822 ( .o(n6310), .a(n6309) );
no02f01  g0823 ( .o(n6311_1), .a(n6310), .b(_net_274) );
no02f01  g0824 ( .o(n6312), .a(n6309), .b(n5522) );
oa12f01  g0825 ( .o(n6313), .a(n6190), .b(n6312), .c(n6311_1) );
na02f01  g0826 ( .o(n6314), .a(n6207), .b(_net_274) );
na02f01  g0827 ( .o(n6315), .a(n6314), .b(n6313) );
na02f01  g0828 ( .o(n6316_1), .a(n6315), .b(n6308) );
na03f01  g0829 ( .o(n6317), .a(n6314), .b(n6313), .c(net_9431) );
na04f01  g0830 ( .o(n6318), .a(n6317), .b(n6316_1), .c(n6307), .d(n6297_1) );
na02f01  g0831 ( .o(n6319), .a(n6309), .b(_net_274) );
no02f01  g0832 ( .o(n6320), .a(n6319), .b(_net_275) );
ao12f01  g0833 ( .o(n6321_1), .a(n5534), .b(n6309), .c(_net_274) );
oa12f01  g0834 ( .o(n6322), .a(n6190), .b(n6321_1), .c(n6320) );
na02f01  g0835 ( .o(n6323), .a(n6207), .b(_net_275) );
na03f01  g0836 ( .o(n6324), .a(n6323), .b(n6322), .c(net_9432) );
in01f01  g0837 ( .o(n6325), .a(net_9432) );
na02f01  g0838 ( .o(n6326_1), .a(n6323), .b(n6322) );
na02f01  g0839 ( .o(n6327), .a(n6326_1), .b(n6325) );
na02f01  g0840 ( .o(n6328), .a(n6327), .b(n6324) );
in01f01  g0841 ( .o(n6329), .a(net_9433) );
na02f01  g0842 ( .o(n6330), .a(n6207), .b(_net_276) );
no03f01  g0843 ( .o(n6331_1), .a(n6319), .b(_net_276), .c(n5534) );
no02f01  g0844 ( .o(n6332), .a(n6319), .b(n5534) );
no02f01  g0845 ( .o(n6333), .a(n6332), .b(n5579) );
oa12f01  g0846 ( .o(n6334), .a(n6190), .b(n6333), .c(n6331_1) );
ao12f01  g0847 ( .o(n6335), .a(n6329), .b(n6334), .c(n6330) );
na02f01  g0848 ( .o(n6336_1), .a(n6334), .b(n6330) );
no02f01  g0849 ( .o(n6337), .a(n6336_1), .b(net_9433) );
in01f01  g0850 ( .o(n6338), .a(net_9436) );
na02f01  g0851 ( .o(n6339), .a(n6207), .b(net_279) );
no02f01  g0852 ( .o(n6340), .a(n6215), .b(n5543) );
no02f01  g0853 ( .o(n6341_1), .a(n6340), .b(n5594_1) );
no03f01  g0854 ( .o(n6342), .a(n6215), .b(net_279), .c(n5543) );
oa12f01  g0855 ( .o(n6343), .a(n6190), .b(n6342), .c(n6341_1) );
ao12f01  g0856 ( .o(n6344), .a(n6338), .b(n6343), .c(n6339) );
na02f01  g0857 ( .o(n6345), .a(n6343), .b(n6339) );
no02f01  g0858 ( .o(n6346_1), .a(n6345), .b(net_9436) );
oa22f01  g0859 ( .o(n6347), .a(n6346_1), .b(n6344), .c(n6337), .d(n6335) );
no04f01  g0860 ( .o(n6348), .a(n6347), .b(n6328), .c(n6318), .d(n6224) );
no02f01  g0861 ( .o(n6349), .a(net_9539), .b(net_9513) );
na02f01  g0862 ( .o(n6350), .a(n6349), .b(n6221_1) );
in01f01  g0863 ( .o(n6351_1), .a(n6349) );
na02f01  g0864 ( .o(n6352), .a(n6351_1), .b(_net_9266) );
oa12f01  g0865 ( .o(n613), .a(n6352), .b(n6350), .c(n6348) );
in01f01  g0866 ( .o(n6354), .a(net_9310) );
in01f01  g0867 ( .o(n6355), .a(_net_9302) );
no02f01  g0868 ( .o(n6356_1), .a(_net_9301), .b(n6355) );
in01f01  g0869 ( .o(n6357), .a(_net_9301) );
no02f01  g0870 ( .o(n6358), .a(n6357), .b(_net_9302) );
no02f01  g0871 ( .o(n6359), .a(n6358), .b(n6356_1) );
in01f01  g0872 ( .o(n6360_1), .a(n6359) );
no02f01  g0873 ( .o(n6361), .a(n6360_1), .b(net_9303) );
in01f01  g0874 ( .o(n6362), .a(net_9303) );
no02f01  g0875 ( .o(n6363), .a(n6359), .b(n6362) );
no02f01  g0876 ( .o(n6364_1), .a(n6363), .b(n6361) );
in01f01  g0877 ( .o(n6365), .a(n6364_1) );
no02f01  g0878 ( .o(n6366), .a(n6365), .b(net_9304) );
in01f01  g0879 ( .o(n6367), .a(net_9304) );
no02f01  g0880 ( .o(n6368), .a(n6364_1), .b(n6367) );
no02f01  g0881 ( .o(n6369_1), .a(n6368), .b(n6366) );
in01f01  g0882 ( .o(n6370), .a(n6369_1) );
no02f01  g0883 ( .o(n6371), .a(net_195), .b(n5783) );
no02f01  g0884 ( .o(n6372), .a(n5787_1), .b(_net_193) );
in01f01  g0885 ( .o(n6373_1), .a(net_9307) );
no02f01  g0886 ( .o(n6374), .a(n6373_1), .b(net_9358) );
na02f01  g0887 ( .o(n6375), .a(n6373_1), .b(net_9358) );
in01f01  g0888 ( .o(n6376), .a(n6375) );
no04f01  g0889 ( .o(n6377), .a(n6376), .b(n6374), .c(n6372), .d(n6371) );
no02f01  g0890 ( .o(n6378_1), .a(n6372), .b(n6371) );
in01f01  g0891 ( .o(n6379), .a(n6374) );
ao12f01  g0892 ( .o(n6380), .a(n6378_1), .b(n6375), .c(n6379) );
no02f01  g0893 ( .o(n6381), .a(n6380), .b(n6377) );
in01f01  g0894 ( .o(n6382), .a(n6381) );
no02f01  g0895 ( .o(n6383_1), .a(n6382), .b(n6370) );
no02f01  g0896 ( .o(n6384), .a(n6381), .b(n6369_1) );
no02f01  g0897 ( .o(n6385), .a(n6384), .b(n6383_1) );
no02f01  g0898 ( .o(n6386), .a(n5783), .b(net_9305) );
in01f01  g0899 ( .o(n6387), .a(net_9305) );
no02f01  g0900 ( .o(n6388_1), .a(_net_193), .b(n6387) );
no02f01  g0901 ( .o(n6389), .a(n6388_1), .b(n6386) );
in01f01  g0902 ( .o(n6390), .a(n6389) );
no02f01  g0903 ( .o(n6391), .a(net_194), .b(n5791) );
no02f01  g0904 ( .o(n6392), .a(n5779), .b(net_196) );
no02f01  g0905 ( .o(n6393_1), .a(n6392), .b(n6391) );
in01f01  g0906 ( .o(n6394), .a(n6393_1) );
no02f01  g0907 ( .o(n6395), .a(n6394), .b(net_9359) );
na02f01  g0908 ( .o(n6396), .a(n6394), .b(net_9359) );
in01f01  g0909 ( .o(n6397_1), .a(n6396) );
no03f01  g0910 ( .o(n6398), .a(n6397_1), .b(n6395), .c(n6390) );
in01f01  g0911 ( .o(n6399), .a(n6395) );
ao12f01  g0912 ( .o(n6400), .a(n6389), .b(n6396), .c(n6399) );
no02f01  g0913 ( .o(n6401_1), .a(n6400), .b(n6398) );
in01f01  g0914 ( .o(n6402), .a(n6401_1) );
no02f01  g0915 ( .o(n6403), .a(n6402), .b(n6370) );
no02f01  g0916 ( .o(n6404), .a(n6401_1), .b(n6369_1) );
no02f01  g0917 ( .o(n6405), .a(n6373_1), .b(net_194) );
no02f01  g0918 ( .o(n6406_1), .a(net_9307), .b(n5779) );
in01f01  g0919 ( .o(n6407), .a(net_9306) );
no02f01  g0920 ( .o(n6408), .a(n6407), .b(net_9357) );
na02f01  g0921 ( .o(n6409), .a(n6407), .b(net_9357) );
in01f01  g0922 ( .o(n6410), .a(n6409) );
no04f01  g0923 ( .o(n6411_1), .a(n6410), .b(n6408), .c(n6406_1), .d(n6405) );
no02f01  g0924 ( .o(n6412), .a(n6406_1), .b(n6405) );
in01f01  g0925 ( .o(n6413), .a(n6408) );
ao12f01  g0926 ( .o(n6414), .a(n6412), .b(n6409), .c(n6413) );
no02f01  g0927 ( .o(n6415), .a(n6414), .b(n6411_1) );
in01f01  g0928 ( .o(n6416_1), .a(n6415) );
no02f01  g0929 ( .o(n6417), .a(n6416_1), .b(n6365) );
no02f01  g0930 ( .o(n6418), .a(n6415), .b(n6364_1) );
no02f01  g0931 ( .o(n6419), .a(n6418), .b(n6417) );
no02f01  g0932 ( .o(n6420), .a(n6373_1), .b(net_9305) );
no02f01  g0933 ( .o(n6421_1), .a(net_9307), .b(n6387) );
no02f01  g0934 ( .o(n6422), .a(_net_9301), .b(n6367) );
no02f01  g0935 ( .o(n6423), .a(n6357), .b(net_9304) );
no04f01  g0936 ( .o(n6424), .a(n6423), .b(n6422), .c(n6421_1), .d(n6420) );
no02f01  g0937 ( .o(n6425), .a(n6421_1), .b(n6420) );
no02f01  g0938 ( .o(n6426_1), .a(n6423), .b(n6422) );
no02f01  g0939 ( .o(n6427), .a(n6426_1), .b(n6425) );
no02f01  g0940 ( .o(n6428), .a(net_195), .b(net_9360) );
na02f01  g0941 ( .o(n6429), .a(net_195), .b(net_9360) );
in01f01  g0942 ( .o(n6430), .a(n6429) );
no02f01  g0943 ( .o(n6431_1), .a(n6430), .b(n6428) );
in01f01  g0944 ( .o(n6432), .a(n6431_1) );
no03f01  g0945 ( .o(n6433), .a(n6432), .b(n6427), .c(n6424) );
no02f01  g0946 ( .o(n6434), .a(n6427), .b(n6424) );
no02f01  g0947 ( .o(n6435), .a(n6431_1), .b(n6434) );
no02f01  g0948 ( .o(n6436_1), .a(n6435), .b(n6433) );
no02f01  g0949 ( .o(n6437), .a(net_9361), .b(net_196) );
na02f01  g0950 ( .o(n6438), .a(net_9361), .b(net_196) );
in01f01  g0951 ( .o(n6439), .a(n6438) );
no03f01  g0952 ( .o(n6440), .a(n6439), .b(n6437), .c(net_9306) );
in01f01  g0953 ( .o(n6441_1), .a(n6437) );
ao12f01  g0954 ( .o(n6442), .a(n6407), .b(n6438), .c(n6441_1) );
no02f01  g0955 ( .o(n6443), .a(n6442), .b(n6440) );
no02f01  g0956 ( .o(n6444), .a(n6390), .b(n6360_1) );
no02f01  g0957 ( .o(n6445), .a(n6389), .b(n6359) );
no02f01  g0958 ( .o(n6446_1), .a(n6445), .b(n6444) );
no02f01  g0959 ( .o(n6447), .a(n6446_1), .b(n6443) );
na02f01  g0960 ( .o(n6448), .a(n6446_1), .b(n6443) );
in01f01  g0961 ( .o(n6449), .a(n6448) );
no04f01  g0962 ( .o(n6450), .a(n6449), .b(n6447), .c(n6436_1), .d(n6419) );
oa12f01  g0963 ( .o(n6451_1), .a(n6450), .b(n6404), .c(n6403) );
no02f01  g0964 ( .o(n6452), .a(n6451_1), .b(n6385) );
no02f01  g0965 ( .o(n5633), .a(n6452), .b(n6354) );
in01f01  g0966 ( .o(n6454), .a(_net_9343) );
no02f01  g0967 ( .o(n6455), .a(n6454), .b(_net_9344) );
in01f01  g0968 ( .o(n6456_1), .a(n6455) );
in01f01  g0969 ( .o(n6457), .a(_net_9345) );
no02f01  g0970 ( .o(n6458), .a(n6457), .b(_net_9346) );
in01f01  g0971 ( .o(n6459), .a(n6458) );
no02f01  g0972 ( .o(n6460_1), .a(n6459), .b(n6456_1) );
in01f01  g0973 ( .o(n6461), .a(n6460_1) );
no03f01  g0974 ( .o(n618), .a(n6461), .b(n5633), .c(n6354) );
in01f01  g0975 ( .o(n6463), .a(_net_9238) );
na02f01  g0976 ( .o(n6464_1), .a(net_9233), .b(_net_9167) );
in01f01  g0977 ( .o(n6465), .a(_net_9196) );
no02f01  g0978 ( .o(n1774), .a(n6465), .b(_net_9195) );
na02f01  g0979 ( .o(n6467), .a(n1774), .b(net_9199) );
in01f01  g0980 ( .o(n6468), .a(n6467) );
in01f01  g0981 ( .o(n6469_1), .a(_net_9165) );
no02f01  g0982 ( .o(n6136), .a(_net_9196), .b(_net_9195) );
na02f01  g0983 ( .o(n6471), .a(n6136), .b(net_9200) );
no02f01  g0984 ( .o(n6472), .a(n6471), .b(n6469_1) );
no02f01  g0985 ( .o(n6473), .a(n6472), .b(n6468) );
na02f01  g0986 ( .o(n6474_1), .a(n6473), .b(n6464_1) );
in01f01  g0987 ( .o(n6475), .a(_net_9245) );
no02f01  g0988 ( .o(n6476), .a(net_9170), .b(n6475) );
in01f01  g0989 ( .o(n6477), .a(n6476) );
ao12f01  g0990 ( .o(n6478), .a(n6463), .b(n6477), .c(n6474_1) );
in01f01  g0991 ( .o(n6479_1), .a(_net_9237) );
in01f01  g0992 ( .o(n6480), .a(_net_9171) );
in01f01  g0993 ( .o(n6481), .a(_net_9195) );
no02f01  g0994 ( .o(n7489), .a(_net_9196), .b(n6481) );
na02f01  g0995 ( .o(n6483), .a(n7489), .b(net_9198) );
no02f01  g0996 ( .o(n6484_1), .a(n6483), .b(n6480) );
no02f01  g0997 ( .o(n6485), .a(n6471), .b(n6480) );
in01f01  g0998 ( .o(n6486), .a(n6485) );
oa12f01  g0999 ( .o(n6487), .a(n6486), .b(n6484_1), .c(_net_9238) );
no02f01  g1000 ( .o(n6488), .a(n6487), .b(n6479_1) );
in01f01  g1001 ( .o(n6489_1), .a(_net_9241) );
no02f01  g1002 ( .o(n6490), .a(n6489_1), .b(_net_9171) );
in01f01  g1003 ( .o(n6491), .a(_net_9239) );
no02f01  g1004 ( .o(n6492), .a(n6136), .b(n6491) );
no02f01  g1005 ( .o(n6493_1), .a(n6492), .b(n6490) );
in01f01  g1006 ( .o(n6494), .a(n6493_1) );
in01f01  g1007 ( .o(n6495), .a(_net_9240) );
no02f01  g1008 ( .o(n6496), .a(n6495), .b(_net_9172) );
no02f01  g1009 ( .o(n6497), .a(_net_9244), .b(_net_9242) );
no02f01  g1010 ( .o(n6498_1), .a(n6497), .b(_net_9169) );
no02f01  g1011 ( .o(n6499), .a(n6498_1), .b(n6496) );
in01f01  g1012 ( .o(n6500), .a(n6499) );
oa12f01  g1013 ( .o(n6501), .a(_net_9238), .b(n6500), .c(n6494) );
in01f01  g1014 ( .o(n6502), .a(n6471) );
no02f01  g1015 ( .o(n6503_1), .a(n6502), .b(n6463) );
in01f01  g1016 ( .o(n6504), .a(_net_9247) );
in01f01  g1017 ( .o(n6505), .a(n6483) );
no03f01  g1018 ( .o(n6506), .a(n6505), .b(_net_9176), .c(n6504) );
in01f01  g1019 ( .o(n6507_1), .a(_net_9246) );
no03f01  g1020 ( .o(n6508), .a(n6468), .b(_net_9176), .c(n6507_1) );
oa12f01  g1021 ( .o(n6509), .a(n6503_1), .b(n6508), .c(n6506) );
na02f01  g1022 ( .o(n6510), .a(n6509), .b(n6501) );
in01f01  g1023 ( .o(n6511), .a(_net_9236) );
in01f01  g1024 ( .o(n6512_1), .a(_net_9166) );
no02f01  g1025 ( .o(n6513), .a(n6512_1), .b(net_313) );
in01f01  g1026 ( .o(n6514), .a(net_313) );
in01f01  g1027 ( .o(n6515), .a(_net_9194) );
na04f01  g1028 ( .o(n6516), .a(_net_9165), .b(_net_9168), .c(n6515), .d(n6514) );
no02f01  g1029 ( .o(n6517_1), .a(n6512_1), .b(n6514) );
no02f01  g1030 ( .o(n6518), .a(n6517_1), .b(n6463) );
oa12f01  g1031 ( .o(n6519), .a(n6516), .b(n6518), .c(n6513) );
in01f01  g1032 ( .o(n6520), .a(_net_9243) );
no03f01  g1033 ( .o(n6521), .a(_net_9209), .b(n6520), .c(n6463) );
ao12f01  g1034 ( .o(n6522_1), .a(n6521), .b(n6503_1), .c(_net_9248) );
oa12f01  g1035 ( .o(n6523), .a(n6522_1), .b(n6519), .c(n6511) );
no04f01  g1036 ( .o(n6524), .a(n6523), .b(n6510), .c(n6488), .d(n6478) );
no02f01  g1037 ( .o(n6525), .a(x3390), .b(n5658) );
in01f01  g1038 ( .o(n6526_1), .a(n6525) );
no02f01  g1039 ( .o(n623), .a(n6526_1), .b(n6524) );
no02f01  g1040 ( .o(n6528), .a(n5903_1), .b(n5660) );
in01f01  g1041 ( .o(n6529), .a(net_10490) );
no02f01  g1042 ( .o(n6530), .a(n5675), .b(n6529) );
in01f01  g1043 ( .o(n6531_1), .a(n6530) );
no03f01  g1044 ( .o(n6532), .a(n6531_1), .b(n6528), .c(n5658) );
ao12f01  g1045 ( .o(n6533), .a(n5658), .b(n6532), .c(net_247) );
no03f01  g1046 ( .o(n6534), .a(n6530), .b(n6528), .c(n5658) );
no03f01  g1047 ( .o(n6535), .a(n5903_1), .b(n5660), .c(n5658) );
ao22f01  g1048 ( .o(n6536_1), .a(n6535), .b(x5077), .c(n6534), .d(net_10007) );
na02f01  g1049 ( .o(n633), .a(n6536_1), .b(n6533) );
in01f01  g1050 ( .o(n6538), .a(net_9619) );
in01f01  g1051 ( .o(n6539), .a(net_9618) );
in01f01  g1052 ( .o(n6540), .a(net_9617) );
in01f01  g1053 ( .o(n6541_1), .a(net_9614) );
in01f01  g1054 ( .o(n6542), .a(net_9615) );
no02f01  g1055 ( .o(n6543), .a(n6542), .b(n6541_1) );
na02f01  g1056 ( .o(n6544), .a(n6543), .b(net_9616) );
no02f01  g1057 ( .o(n6545), .a(n6544), .b(n6540) );
in01f01  g1058 ( .o(n6546_1), .a(n6545) );
no02f01  g1059 ( .o(n6547), .a(n6546_1), .b(n6539) );
in01f01  g1060 ( .o(n6548), .a(n6547) );
no02f01  g1061 ( .o(n6549), .a(n6548), .b(n6538) );
in01f01  g1062 ( .o(n6550), .a(net_9613) );
oa12f01  g1063 ( .o(n6551_1), .a(n6550), .b(n6547), .c(net_9619) );
no02f01  g1064 ( .o(n642), .a(n6551_1), .b(n6549) );
no03f01  g1065 ( .o(n6553), .a(n5899), .b(n5631), .c(x6351) );
in01f01  g1066 ( .o(n6554), .a(n6553) );
no02f01  g1067 ( .o(n6555), .a(n6554), .b(n5771) );
in01f01  g1068 ( .o(n6556_1), .a(net_10081) );
in01f01  g1069 ( .o(n6557), .a(net_209) );
no03f01  g1070 ( .o(n6558), .a(n5666_1), .b(x6401), .c(x6445) );
in01f01  g1071 ( .o(n6559), .a(n6558) );
no02f01  g1072 ( .o(n6560), .a(n5549), .b(x6577) );
in01f01  g1073 ( .o(n6561_1), .a(n6560) );
no02f01  g1074 ( .o(n6562), .a(n6561_1), .b(n6559) );
in01f01  g1075 ( .o(n6563), .a(n6562) );
no02f01  g1076 ( .o(n6564), .a(n6559), .b(n5771) );
in01f01  g1077 ( .o(n6565), .a(n6564) );
oa22f01  g1078 ( .o(n6566_1), .a(n6565), .b(n6556_1), .c(n6563), .d(n6557) );
ao12f01  g1079 ( .o(n6567), .a(n6566_1), .b(n6555), .c(net_9975) );
no04f01  g1080 ( .o(n6568), .a(x6496), .b(n5564), .c(n5631), .d(x6351) );
in01f01  g1081 ( .o(n6569), .a(n6568) );
no02f01  g1082 ( .o(n6570), .a(x6531), .b(n5655) );
in01f01  g1083 ( .o(n6571_1), .a(n6570) );
no02f01  g1084 ( .o(n6572), .a(n6571_1), .b(n6569) );
no02f01  g1085 ( .o(n6573), .a(n6569), .b(n5771) );
ao22f01  g1086 ( .o(n6574), .a(n6573), .b(net_9876), .c(n6572), .d(net_10392) );
no04f01  g1087 ( .o(n6575_1), .a(x6496), .b(n5564), .c(x6445), .d(x6351) );
in01f01  g1088 ( .o(n6576), .a(n6575_1) );
no02f01  g1089 ( .o(n6577), .a(n6576), .b(n5771) );
no03f01  g1090 ( .o(n6578), .a(n5899), .b(x6445), .c(x6351) );
in01f01  g1091 ( .o(n6579_1), .a(n6578) );
no02f01  g1092 ( .o(n6580), .a(n6579_1), .b(n5660) );
ao22f01  g1093 ( .o(n6581), .a(n6580), .b(net_9809), .c(n6577), .d(net_9678) );
no02f01  g1094 ( .o(n6582), .a(n6569), .b(n5660) );
na02f01  g1095 ( .o(n6583), .a(n6582), .b(net_9908) );
no02f01  g1096 ( .o(n6584_1), .a(n6579_1), .b(n5771) );
no02f01  g1097 ( .o(n6585), .a(n6576), .b(n5660) );
ao22f01  g1098 ( .o(n6586), .a(n6585), .b(net_9710), .c(n6584_1), .d(net_9777) );
na02f01  g1099 ( .o(n6587), .a(n6586), .b(n6583) );
in01f01  g1100 ( .o(n6588), .a(net_10038) );
in01f01  g1101 ( .o(n6589_1), .a(net_10182) );
no02f01  g1102 ( .o(n6590), .a(n6554), .b(n5686) );
in01f01  g1103 ( .o(n6591), .a(n6590) );
no02f01  g1104 ( .o(n6592), .a(n6576), .b(n6571_1) );
in01f01  g1105 ( .o(n6593), .a(n6592) );
oa22f01  g1106 ( .o(n6594_1), .a(n6593), .b(n6589_1), .c(n6591), .d(n6588) );
in01f01  g1107 ( .o(n6595), .a(net_9840) );
in01f01  g1108 ( .o(n6596), .a(net_9741) );
no02f01  g1109 ( .o(n6597), .a(n6576), .b(n5686) );
in01f01  g1110 ( .o(n6598), .a(n6597) );
no02f01  g1111 ( .o(n6599_1), .a(n6579_1), .b(n5686) );
in01f01  g1112 ( .o(n6600), .a(n6599_1) );
oa22f01  g1113 ( .o(n6601), .a(n6600), .b(n6595), .c(n6598), .d(n6596) );
no02f01  g1114 ( .o(n6602), .a(n6554), .b(n5660) );
no02f01  g1115 ( .o(n6603), .a(n6571_1), .b(n6554) );
ao22f01  g1116 ( .o(n6604_1), .a(n6603), .b(net_10497), .c(n6602), .d(net_10007) );
no02f01  g1117 ( .o(n6605), .a(n6579_1), .b(n6571_1) );
no02f01  g1118 ( .o(n6606), .a(n6569), .b(n5686) );
ao22f01  g1119 ( .o(n6607), .a(n6606), .b(net_9939), .c(n6605), .d(net_10287) );
na02f01  g1120 ( .o(n6608), .a(n6607), .b(n6604_1) );
no04f01  g1121 ( .o(n6609_1), .a(n6608), .b(n6601), .c(n6594_1), .d(n6587) );
na04f01  g1122 ( .o(n647), .a(n6609_1), .b(n6581), .c(n6574), .d(n6567) );
no02f01  g1123 ( .o(n6611), .a(n5997), .b(net_9596) );
in01f01  g1124 ( .o(n6612), .a(n6611) );
in01f01  g1125 ( .o(n6613), .a(net_9595) );
in01f01  g1126 ( .o(n6614_1), .a(n5958) );
no02f01  g1127 ( .o(n6615), .a(n6614_1), .b(n6613) );
in01f01  g1128 ( .o(n6616), .a(net_9592) );
in01f01  g1129 ( .o(n6617), .a(n5965) );
no02f01  g1130 ( .o(n6618), .a(n6617), .b(n6616) );
na02f01  g1131 ( .o(n6619_1), .a(n5941), .b(_net_9591) );
no02f01  g1132 ( .o(n6620), .a(n5938), .b(_net_9590) );
no02f01  g1133 ( .o(n6621), .a(n5941), .b(_net_9591) );
no02f01  g1134 ( .o(n6622), .a(n6621), .b(n6620) );
ao12f01  g1135 ( .o(n6623), .a(n6622), .b(n5941), .c(_net_9591) );
in01f01  g1136 ( .o(n6624_1), .a(_net_9590) );
in01f01  g1137 ( .o(n6625), .a(n5938) );
no02f01  g1138 ( .o(n6626), .a(n6625), .b(n6624_1) );
no02f01  g1139 ( .o(n6627), .a(n5945), .b(_net_9589) );
na02f01  g1140 ( .o(n6628), .a(n5945), .b(_net_9589) );
na02f01  g1141 ( .o(n6629_1), .a(n5948), .b(_net_9588) );
ao12f01  g1142 ( .o(n6630), .a(n6627), .b(n6629_1), .c(n6628) );
no02f01  g1143 ( .o(n6631), .a(n6630), .b(n6626) );
ao12f01  g1144 ( .o(n6632), .a(n6623), .b(n6631), .c(n6619_1) );
in01f01  g1145 ( .o(n6633), .a(net_9594) );
in01f01  g1146 ( .o(n6634_1), .a(n5961) );
no02f01  g1147 ( .o(n6635), .a(n6634_1), .b(n6633) );
na02f01  g1148 ( .o(n6636), .a(n5968), .b(net_9593) );
in01f01  g1149 ( .o(n6637), .a(n6636) );
no04f01  g1150 ( .o(n6638), .a(n6637), .b(n6635), .c(n6632), .d(n6618) );
no02f01  g1151 ( .o(n6639_1), .a(n5968), .b(net_9593) );
no02f01  g1152 ( .o(n6640), .a(n5965), .b(net_9592) );
ao12f01  g1153 ( .o(n6641), .a(n6639_1), .b(n6640), .c(n6636) );
no02f01  g1154 ( .o(n6642), .a(n6641), .b(n6635) );
no02f01  g1155 ( .o(n6643), .a(n5961), .b(net_9594) );
no02f01  g1156 ( .o(n6644_1), .a(n5958), .b(net_9595) );
no02f01  g1157 ( .o(n6645), .a(n6644_1), .b(n6643) );
ao12f01  g1158 ( .o(n6646), .a(n6645), .b(n6615), .c(net_9595) );
no02f01  g1159 ( .o(n6647), .a(n6646), .b(n6642) );
in01f01  g1160 ( .o(n6648), .a(n6647) );
no02f01  g1161 ( .o(n6649_1), .a(n6648), .b(n6638) );
no02f01  g1162 ( .o(n6650), .a(n6649_1), .b(n6615) );
na02f01  g1163 ( .o(n6651), .a(n6646), .b(n6614_1) );
in01f01  g1164 ( .o(n6652), .a(n6651) );
no02f01  g1165 ( .o(n6653), .a(n6652), .b(n6650) );
na02f01  g1166 ( .o(n6654_1), .a(n5997), .b(net_9596) );
in01f01  g1167 ( .o(n6655), .a(n6654_1) );
oa12f01  g1168 ( .o(n6656), .a(n6612), .b(n6655), .c(n6653) );
in01f01  g1169 ( .o(n6657), .a(net_9597) );
no02f01  g1170 ( .o(n6658), .a(n5994), .b(n6657) );
no02f01  g1171 ( .o(n6659_1), .a(n5993_1), .b(net_9597) );
no02f01  g1172 ( .o(n6660), .a(n6659_1), .b(n6658) );
in01f01  g1173 ( .o(n6661), .a(n6660) );
na02f01  g1174 ( .o(n6662), .a(n6661), .b(n6656) );
in01f01  g1175 ( .o(n6663), .a(n6653) );
na02f01  g1176 ( .o(n6664_1), .a(n6654_1), .b(n6663) );
na03f01  g1177 ( .o(n6665), .a(n6660), .b(n6664_1), .c(n6612) );
na02f01  g1178 ( .o(n652), .a(n6665), .b(n6662) );
in01f01  g1179 ( .o(n6667), .a(_net_10125) );
na02f01  g1180 ( .o(n6668), .a(n5762), .b(n6667) );
na02f01  g1181 ( .o(n6669_1), .a(n5763_1), .b(_net_10125) );
na02f01  g1182 ( .o(n661), .a(n6669_1), .b(n6668) );
in01f01  g1183 ( .o(n6671), .a(net_9206) );
in01f01  g1184 ( .o(n6672), .a(net_9218) );
in01f01  g1185 ( .o(n6673), .a(n6516) );
no02f01  g1186 ( .o(n6674_1), .a(n6512_1), .b(n6514) );
oa12f01  g1187 ( .o(n6675), .a(_net_9236), .b(n6674_1), .c(n6673) );
na02f01  g1188 ( .o(n6676), .a(n6136), .b(_net_9239) );
in01f01  g1189 ( .o(n6677), .a(_net_9172) );
no02f01  g1190 ( .o(n6678), .a(n6495), .b(n6677) );
in01f01  g1191 ( .o(n6679_1), .a(n6678) );
ao12f01  g1192 ( .o(n6680), .a(_net_9235), .b(_net_9244), .c(_net_9169) );
na04f01  g1193 ( .o(n6681), .a(n6680), .b(n6679_1), .c(n6676), .d(n6675) );
na02f01  g1194 ( .o(n6682), .a(n6472), .b(_net_9238) );
oa12f01  g1195 ( .o(n6683), .a(n6682), .b(n6486), .c(n6479_1) );
no02f01  g1196 ( .o(n6684_1), .a(n6683), .b(n6681) );
oa12f01  g1197 ( .o(n6685), .a(n6684_1), .b(_net_9209), .c(n6672) );
in01f01  g1198 ( .o(n6686), .a(n6684_1) );
no03f01  g1199 ( .o(n6687), .a(n6686), .b(_net_9209), .c(n6672) );
in01f01  g1200 ( .o(n6688), .a(n6687) );
in01f01  g1201 ( .o(n6689_1), .a(net_9205) );
in01f01  g1202 ( .o(n6690), .a(_net_9204) );
in01f01  g1203 ( .o(n6691), .a(_net_9203) );
in01f01  g1204 ( .o(n6692), .a(_net_9202) );
in01f01  g1205 ( .o(n6693), .a(_net_9201) );
no02f01  g1206 ( .o(n6694_1), .a(n6693), .b(n6692) );
in01f01  g1207 ( .o(n6695), .a(n6694_1) );
no02f01  g1208 ( .o(n6696), .a(n6695), .b(n6691) );
in01f01  g1209 ( .o(n6697), .a(n6696) );
no02f01  g1210 ( .o(n6698), .a(n6697), .b(n6690) );
in01f01  g1211 ( .o(n6699_1), .a(n6698) );
no02f01  g1212 ( .o(n6700), .a(n6699_1), .b(n6689_1) );
in01f01  g1213 ( .o(n6701), .a(n6700) );
na02f01  g1214 ( .o(n6702), .a(n6701), .b(n6671) );
no02f01  g1215 ( .o(n6703), .a(n6701), .b(n6671) );
in01f01  g1216 ( .o(n6704_1), .a(n6703) );
na02f01  g1217 ( .o(n6705), .a(n6704_1), .b(n6702) );
oa22f01  g1218 ( .o(n666), .a(n6705), .b(n6688), .c(n6685), .d(n6671) );
in01f01  g1219 ( .o(n6707), .a(_net_10110) );
ao12f01  g1220 ( .o(n6708), .a(n5658), .b(n6160_1), .c(x5143) );
oa12f01  g1221 ( .o(n671), .a(n6708), .b(n6159), .c(n6707) );
in01f01  g1222 ( .o(n1032), .a(_net_10429) );
ao12f01  g1223 ( .o(n6711), .a(n5658), .b(n6052_1), .c(x4851) );
oa12f01  g1224 ( .o(n676), .a(n6711), .b(n6048), .c(n1032) );
in01f01  g1225 ( .o(n6713_1), .a(_net_10143) );
in01f01  g1226 ( .o(n6714), .a(_net_10142) );
no02f01  g1227 ( .o(n6715), .a(n6714), .b(_net_9730) );
in01f01  g1228 ( .o(n6716), .a(n6715) );
oa12f01  g1229 ( .o(n6717), .a(n6713_1), .b(n6716), .c(_net_9731) );
oa12f01  g1230 ( .o(n6718_1), .a(_net_9731), .b(n6716), .c(n6713_1) );
na02f01  g1231 ( .o(n6719), .a(n6718_1), .b(n6717) );
in01f01  g1232 ( .o(n6720), .a(_net_9731) );
no02f01  g1233 ( .o(n6721), .a(_net_10143), .b(n6720) );
in01f01  g1234 ( .o(n6722), .a(n6721) );
in01f01  g1235 ( .o(n6723_1), .a(_net_9730) );
no02f01  g1236 ( .o(n6724), .a(_net_10142), .b(n6723_1) );
in01f01  g1237 ( .o(n6725), .a(_net_10141) );
no02f01  g1238 ( .o(n6726), .a(n6725), .b(_net_9729) );
in01f01  g1239 ( .o(n6727), .a(_net_9728) );
no02f01  g1240 ( .o(n6728_1), .a(_net_10140), .b(n6727) );
in01f01  g1241 ( .o(n6729), .a(_net_9729) );
no02f01  g1242 ( .o(n6730), .a(_net_10141), .b(n6729) );
no02f01  g1243 ( .o(n6731), .a(n6730), .b(n6728_1) );
no02f01  g1244 ( .o(n6732), .a(n6731), .b(n6726) );
no02f01  g1245 ( .o(n6733_1), .a(n6732), .b(n6724) );
na02f01  g1246 ( .o(n6734), .a(n6733_1), .b(n6722) );
na02f01  g1247 ( .o(n6735), .a(n6734), .b(n6719) );
in01f01  g1248 ( .o(n6736), .a(_net_9732) );
no02f01  g1249 ( .o(n6737), .a(n6736), .b(_net_10144) );
in01f01  g1250 ( .o(n6738_1), .a(_net_10144) );
no02f01  g1251 ( .o(n6739), .a(_net_9732), .b(n6738_1) );
no02f01  g1252 ( .o(n6740), .a(n6739), .b(n6737) );
in01f01  g1253 ( .o(n6741), .a(net_10199) );
no02f01  g1254 ( .o(n6742), .a(n6031), .b(n5674) );
in01f01  g1255 ( .o(n6743_1), .a(n6742) );
oa12f01  g1256 ( .o(n6744), .a(net_10175), .b(_net_133), .c(net_8832) );
na03f01  g1257 ( .o(n6745), .a(n6744), .b(n6743_1), .c(n6741) );
na03f01  g1258 ( .o(n6746), .a(n6745), .b(_net_9740), .c(n6741) );
ao12f01  g1259 ( .o(n6747), .a(n6746), .b(n6740), .c(n6735) );
oa12f01  g1260 ( .o(n6748_1), .a(n6747), .b(n6740), .c(n6735) );
in01f01  g1261 ( .o(n6749), .a(_net_9740) );
no02f01  g1262 ( .o(n6750), .a(n6749), .b(n6741) );
in01f01  g1263 ( .o(n6751), .a(_net_10140) );
no02f01  g1264 ( .o(n6752), .a(n6751), .b(n6725) );
in01f01  g1265 ( .o(n6753_1), .a(n6752) );
no02f01  g1266 ( .o(n6754), .a(n6753_1), .b(n6714) );
na02f01  g1267 ( .o(n6755), .a(n6754), .b(_net_10143) );
in01f01  g1268 ( .o(n6756), .a(n6755) );
no02f01  g1269 ( .o(n6757), .a(n6756), .b(_net_10144) );
no02f01  g1270 ( .o(n6758_1), .a(n6755), .b(n6738_1) );
no02f01  g1271 ( .o(n6759), .a(n6758_1), .b(n6757) );
no02f01  g1272 ( .o(n6760), .a(n6745), .b(n6749) );
ao22f01  g1273 ( .o(n6761), .a(n6760), .b(_net_10144), .c(n6759), .d(n6750) );
na02f01  g1274 ( .o(n681), .a(n6761), .b(n6748_1) );
no02f01  g1275 ( .o(n6763_1), .a(n6142), .b(n6136_1) );
ao12f01  g1276 ( .o(n6764), .a(n6763_1), .b(n6136_1), .c(_net_9385) );
na04f01  g1277 ( .o(n6765), .a(n6764), .b(n6131_1), .c(_net_9381), .d(x6599) );
in01f01  g1278 ( .o(n6766), .a(n6131_1) );
na04f01  g1279 ( .o(n6767), .a(n6764), .b(n6766), .c(_net_8825), .d(x6599) );
na02f01  g1280 ( .o(n686), .a(n6767), .b(n6765) );
in01f01  g1281 ( .o(n6769), .a(_net_10256) );
in01f01  g1282 ( .o(n6770), .a(_net_10254) );
in01f01  g1283 ( .o(n6771), .a(_net_10253) );
no02f01  g1284 ( .o(n6772), .a(n6771), .b(_net_9835) );
in01f01  g1285 ( .o(n6773_1), .a(_net_9835) );
no02f01  g1286 ( .o(n6774), .a(_net_10253), .b(n6773_1) );
in01f01  g1287 ( .o(n6775), .a(n6774) );
in01f01  g1288 ( .o(n6776), .a(_net_9834) );
no02f01  g1289 ( .o(n6777), .a(_net_10252), .b(n6776) );
in01f01  g1290 ( .o(n6778_1), .a(_net_9831) );
no02f01  g1291 ( .o(n6779), .a(_net_10249), .b(n6778_1) );
in01f01  g1292 ( .o(n6780), .a(_net_10248) );
in01f01  g1293 ( .o(n6781), .a(_net_10247) );
no02f01  g1294 ( .o(n6782_1), .a(_net_9829), .b(n6781) );
no02f01  g1295 ( .o(n6783), .a(_net_9830), .b(n6780) );
no02f01  g1296 ( .o(n6784), .a(n6783), .b(n6782_1) );
in01f01  g1297 ( .o(n6785), .a(_net_9829) );
no02f01  g1298 ( .o(n6786_1), .a(n6785), .b(_net_10247) );
in01f01  g1299 ( .o(n6787), .a(_net_10246) );
no02f01  g1300 ( .o(n6788), .a(n6787), .b(_net_9828) );
no02f01  g1301 ( .o(n6789), .a(_net_10245), .b(n6183) );
no02f01  g1302 ( .o(n6790), .a(_net_10246), .b(n6178) );
no02f01  g1303 ( .o(n6791_1), .a(n6790), .b(n6789) );
no02f01  g1304 ( .o(n6792), .a(n6791_1), .b(n6788) );
no02f01  g1305 ( .o(n6793), .a(n6792), .b(n6786_1) );
in01f01  g1306 ( .o(n6794), .a(n6793) );
ao22f01  g1307 ( .o(n6795), .a(n6794), .b(n6784), .c(_net_9830), .d(n6780) );
in01f01  g1308 ( .o(n6796_1), .a(n6795) );
no02f01  g1309 ( .o(n6797), .a(n6796_1), .b(n6779) );
in01f01  g1310 ( .o(n6798), .a(n6797) );
in01f01  g1311 ( .o(n6799), .a(_net_9833) );
no02f01  g1312 ( .o(n6800), .a(_net_10251), .b(n6799) );
in01f01  g1313 ( .o(n6801_1), .a(_net_9832) );
no02f01  g1314 ( .o(n6802), .a(_net_10250), .b(n6801_1) );
no03f01  g1315 ( .o(n6803), .a(n6802), .b(n6800), .c(n6798) );
in01f01  g1316 ( .o(n6804), .a(n6802) );
in01f01  g1317 ( .o(n6805), .a(_net_10250) );
no02f01  g1318 ( .o(n6806_1), .a(n6805), .b(_net_9832) );
in01f01  g1319 ( .o(n6807), .a(_net_10249) );
no02f01  g1320 ( .o(n6808), .a(n6807), .b(_net_9831) );
ao12f01  g1321 ( .o(n6809), .a(n6806_1), .b(n6808), .c(n6804) );
no02f01  g1322 ( .o(n6810), .a(n6809), .b(n6800) );
in01f01  g1323 ( .o(n6811_1), .a(_net_10251) );
no02f01  g1324 ( .o(n6812), .a(n6811_1), .b(_net_9833) );
in01f01  g1325 ( .o(n6813), .a(_net_10252) );
no02f01  g1326 ( .o(n6814), .a(n6813), .b(_net_9834) );
no02f01  g1327 ( .o(n6815), .a(n6814), .b(n6812) );
ao12f01  g1328 ( .o(n6816_1), .a(n6815), .b(n6777), .c(_net_9834) );
no02f01  g1329 ( .o(n6817), .a(n6816_1), .b(n6810) );
in01f01  g1330 ( .o(n6818), .a(n6817) );
no02f01  g1331 ( .o(n6819), .a(n6818), .b(n6803) );
na02f01  g1332 ( .o(n6820), .a(n6816_1), .b(_net_10252) );
oa12f01  g1333 ( .o(n6821_1), .a(n6820), .b(n6819), .c(n6777) );
ao12f01  g1334 ( .o(n6822), .a(n6772), .b(n6821_1), .c(n6775) );
na02f01  g1335 ( .o(n6823), .a(n6822), .b(n6770) );
no03f01  g1336 ( .o(n6824), .a(n6823), .b(_net_10255), .c(n6769) );
no02f01  g1337 ( .o(n6825), .a(n6823), .b(_net_10255) );
oa12f01  g1338 ( .o(n6826_1), .a(n6177_1), .b(n6825), .c(_net_10256) );
no02f01  g1339 ( .o(n6827), .a(n6805), .b(n6807) );
in01f01  g1340 ( .o(n6828), .a(n6827) );
in01f01  g1341 ( .o(n6829), .a(_net_10245) );
no02f01  g1342 ( .o(n6830), .a(n6787), .b(n6829) );
in01f01  g1343 ( .o(n6831_1), .a(n6830) );
no02f01  g1344 ( .o(n6832), .a(n6831_1), .b(n6781) );
in01f01  g1345 ( .o(n6833), .a(n6832) );
no02f01  g1346 ( .o(n6834), .a(n6833), .b(n6780) );
in01f01  g1347 ( .o(n6835), .a(n6834) );
no02f01  g1348 ( .o(n6836_1), .a(n6835), .b(n6828) );
in01f01  g1349 ( .o(n6837), .a(n6836_1) );
no02f01  g1350 ( .o(n6838), .a(n6837), .b(n6811_1) );
in01f01  g1351 ( .o(n6839), .a(n6838) );
no02f01  g1352 ( .o(n6840), .a(n6839), .b(n6813) );
na02f01  g1353 ( .o(n6841_1), .a(n6840), .b(_net_10253) );
no02f01  g1354 ( .o(n6842), .a(n6841_1), .b(n6770) );
na02f01  g1355 ( .o(n6843), .a(n6842), .b(_net_10255) );
in01f01  g1356 ( .o(n6844), .a(n6843) );
na02f01  g1357 ( .o(n6845), .a(n6844), .b(_net_10256) );
in01f01  g1358 ( .o(n6846_1), .a(n6175) );
ao12f01  g1359 ( .o(n6847), .a(n6846_1), .b(n6843), .c(n6769) );
ao22f01  g1360 ( .o(n6848), .a(n6847), .b(n6845), .c(n6168), .d(_net_10256) );
oa12f01  g1361 ( .o(n691), .a(n6848), .b(n6826_1), .c(n6824) );
no02f01  g1362 ( .o(n6850), .a(n6484_1), .b(n6479_1) );
in01f01  g1363 ( .o(n6851_1), .a(_net_9249) );
no02f01  g1364 ( .o(n6852), .a(n6485), .b(n6851_1) );
in01f01  g1365 ( .o(n6853), .a(_net_9176) );
no02f01  g1366 ( .o(n6854), .a(_net_9176), .b(n6851_1) );
ao22f01  g1367 ( .o(n6855), .a(n6854), .b(n6483), .c(n6502), .d(n6853) );
ao22f01  g1368 ( .o(n6856_1), .a(n6854), .b(n6467), .c(n6502), .d(n6853) );
oa22f01  g1369 ( .o(n6857), .a(n6856_1), .b(n6507_1), .c(n6855), .d(n6504) );
ao12f01  g1370 ( .o(n6858), .a(n6857), .b(n6852), .c(n6850) );
no03f01  g1371 ( .o(n6859), .a(n6474_1), .b(n6851_1), .c(n6463) );
no03f01  g1372 ( .o(n6860), .a(n6517_1), .b(n6673), .c(n6513) );
in01f01  g1373 ( .o(n6861_1), .a(n6860) );
no03f01  g1374 ( .o(n6862), .a(n6861_1), .b(n6511), .c(n6851_1) );
na02f01  g1375 ( .o(n6863), .a(_net_9248), .b(_net_9249) );
in01f01  g1376 ( .o(n6864), .a(_net_9209) );
no02f01  g1377 ( .o(n6865_1), .a(n6520), .b(n6851_1) );
ao22f01  g1378 ( .o(n6866), .a(n6865_1), .b(n6864), .c(n6476), .d(_net_9249) );
oa12f01  g1379 ( .o(n6867), .a(n6866), .b(n6863), .c(n6502) );
ao12f01  g1380 ( .o(n6868), .a(n6851_1), .b(n6499), .c(n6493_1) );
no04f01  g1381 ( .o(n6869), .a(n6868), .b(n6867), .c(n6862), .d(n6859) );
ao12f01  g1382 ( .o(n696), .a(n6526_1), .b(n6869), .c(n6858) );
no02f01  g1383 ( .o(n6871), .a(n5690_1), .b(n5660) );
in01f01  g1384 ( .o(n6872), .a(net_10385) );
no02f01  g1385 ( .o(n6873), .a(n5675), .b(n6872) );
in01f01  g1386 ( .o(n6874), .a(n6873) );
no03f01  g1387 ( .o(n6875_1), .a(n6874), .b(n6871), .c(n5658) );
ao12f01  g1388 ( .o(n6876), .a(n5658), .b(n6875_1), .c(net_260) );
no03f01  g1389 ( .o(n6877), .a(n6873), .b(n6871), .c(n5658) );
no03f01  g1390 ( .o(n6878), .a(n5690_1), .b(n5660), .c(n5658) );
ao22f01  g1391 ( .o(n6879), .a(n6878), .b(x4041), .c(n6877), .d(net_9921) );
na02f01  g1392 ( .o(n701), .a(n6879), .b(n6876) );
in01f01  g1393 ( .o(n3465), .a(_net_10219) );
na04f01  g1394 ( .o(n6882), .a(n5665), .b(x6496), .c(x6401), .d(n5631) );
no02f01  g1395 ( .o(n6883), .a(n6882), .b(n5664) );
no02f01  g1396 ( .o(n6884), .a(n6883), .b(n5658) );
no02f01  g1397 ( .o(n6885_1), .a(n6884), .b(n5768_1) );
in01f01  g1398 ( .o(n6886), .a(n6883) );
no02f01  g1399 ( .o(n6887), .a(n6886), .b(n5773_1) );
ao12f01  g1400 ( .o(n6888), .a(n5658), .b(n6887), .c(x4851) );
oa12f01  g1401 ( .o(n706), .a(n6888), .b(n6885_1), .c(n3465) );
in01f01  g1402 ( .o(n6890_1), .a(net_10034) );
oa22f01  g1403 ( .o(n711), .a(n5907), .b(n6890_1), .c(n5905), .d(n5600) );
na02f01  g1404 ( .o(n6892), .a(n6038), .b(net_238) );
na02f01  g1405 ( .o(n6893), .a(n6037_1), .b(net_9867) );
ao22f01  g1406 ( .o(n6894), .a(n6044), .b(x5647), .c(n6042_1), .d(_net_10312) );
na04f01  g1407 ( .o(n716), .a(n6894), .b(n6893), .c(n6892), .d(n6040) );
ao12f01  g1408 ( .o(n6896), .a(n5658), .b(n6875_1), .c(net_256) );
ao22f01  g1409 ( .o(n6897), .a(n6878), .b(x4359), .c(n6877), .d(net_9917) );
na02f01  g1410 ( .o(n726), .a(n6897), .b(n6896) );
in01f01  g1411 ( .o(n6899), .a(_net_10323) );
ao12f01  g1412 ( .o(n6900_1), .a(n5658), .b(n5774), .c(x4937) );
oa12f01  g1413 ( .o(n731), .a(n6900_1), .b(n5770), .c(n6899) );
in01f01  g1414 ( .o(n6902), .a(_net_10260) );
in01f01  g1415 ( .o(n6903), .a(_net_10259) );
in01f01  g1416 ( .o(n6904), .a(_net_9830) );
oa22f01  g1417 ( .o(n6905_1), .a(n6904), .b(n6902), .c(n6903), .d(n6785) );
no02f01  g1418 ( .o(n6906), .a(_net_10259), .b(_net_9829) );
ao12f01  g1419 ( .o(n6907), .a(n6179), .b(n6184), .c(n6182) );
no02f01  g1420 ( .o(n6908), .a(n6907), .b(n6906) );
oa22f01  g1421 ( .o(n6909), .a(n6908), .b(n6905_1), .c(_net_9830), .d(_net_10260) );
no02f01  g1422 ( .o(n6910_1), .a(_net_10261), .b(_net_9831) );
no02f01  g1423 ( .o(n6911), .a(_net_9833), .b(_net_10263) );
no02f01  g1424 ( .o(n6912), .a(_net_9832), .b(_net_10262) );
no04f01  g1425 ( .o(n6913), .a(n6912), .b(n6911), .c(n6910_1), .d(n6909) );
in01f01  g1426 ( .o(n6914_1), .a(n6911) );
in01f01  g1427 ( .o(n6915), .a(n6912) );
in01f01  g1428 ( .o(n6916), .a(_net_10262) );
no02f01  g1429 ( .o(n6917), .a(n6801_1), .b(n6916) );
in01f01  g1430 ( .o(n6918), .a(_net_10261) );
no02f01  g1431 ( .o(n6919_1), .a(n6918), .b(n6778_1) );
ao12f01  g1432 ( .o(n6920), .a(n6917), .b(n6919_1), .c(n6915) );
in01f01  g1433 ( .o(n6921), .a(n6920) );
na02f01  g1434 ( .o(n6922), .a(n6921), .b(n6914_1) );
in01f01  g1435 ( .o(n6923), .a(_net_10263) );
no02f01  g1436 ( .o(n6924_1), .a(n6799), .b(n6923) );
in01f01  g1437 ( .o(n6925), .a(n6924_1) );
na02f01  g1438 ( .o(n6926), .a(n6925), .b(n6922) );
no02f01  g1439 ( .o(n6927), .a(n6926), .b(n6913) );
in01f01  g1440 ( .o(n6928), .a(_net_10264) );
no02f01  g1441 ( .o(n6929_1), .a(n6776), .b(n6928) );
no02f01  g1442 ( .o(n6930), .a(_net_9834), .b(_net_10264) );
no02f01  g1443 ( .o(n6931), .a(n6930), .b(n6929_1) );
in01f01  g1444 ( .o(n6932), .a(n6931) );
in01f01  g1445 ( .o(n6933), .a(n6177_1) );
ao12f01  g1446 ( .o(n6934_1), .a(n6933), .b(n6932), .c(n6927) );
oa12f01  g1447 ( .o(n6935), .a(n6934_1), .b(n6932), .c(n6927) );
in01f01  g1448 ( .o(n6936), .a(n6170) );
no02f01  g1449 ( .o(n6937), .a(n6936), .b(_net_10259) );
na02f01  g1450 ( .o(n6938), .a(n6937), .b(n6902) );
no02f01  g1451 ( .o(n6939_1), .a(n6938), .b(_net_10261) );
in01f01  g1452 ( .o(n6940), .a(n6939_1) );
no02f01  g1453 ( .o(n6941), .a(n6940), .b(_net_10262) );
in01f01  g1454 ( .o(n6942), .a(n6941) );
no02f01  g1455 ( .o(n6943), .a(n6942), .b(_net_10263) );
in01f01  g1456 ( .o(n6944_1), .a(n6943) );
no02f01  g1457 ( .o(n6945), .a(n6944_1), .b(_net_10264) );
in01f01  g1458 ( .o(n6946), .a(n6945) );
na02f01  g1459 ( .o(n6947), .a(n6944_1), .b(_net_10264) );
na02f01  g1460 ( .o(n6948), .a(n6947), .b(n6946) );
ao22f01  g1461 ( .o(n6949_1), .a(n6948), .b(n6175), .c(n6168), .d(_net_10264) );
na02f01  g1462 ( .o(n741), .a(n6949_1), .b(n6935) );
ao22f01  g1463 ( .o(n6951), .a(n6585), .b(net_9705), .c(n6562), .d(net_208) );
ao22f01  g1464 ( .o(n6952), .a(n6599_1), .b(net_9836), .c(n6584_1), .d(net_9772) );
ao22f01  g1465 ( .o(n6953), .a(n6580), .b(net_9804), .c(n6573), .d(net_9871) );
in01f01  g1466 ( .o(n6954_1), .a(net_9970) );
in01f01  g1467 ( .o(n6955), .a(n6555) );
no02f01  g1468 ( .o(n6956), .a(n6955), .b(n6954_1) );
in01f01  g1469 ( .o(n6957), .a(net_10002) );
in01f01  g1470 ( .o(n6958_1), .a(net_9737) );
in01f01  g1471 ( .o(n6959), .a(n6602) );
oa22f01  g1472 ( .o(n6960), .a(n6959), .b(n6957), .c(n6598), .d(n6958_1) );
na02f01  g1473 ( .o(n6961), .a(n6577), .b(net_9673) );
oa12f01  g1474 ( .o(n6962_1), .a(n6961), .b(n6591), .c(n6890_1) );
in01f01  g1475 ( .o(n6963), .a(net_9903) );
in01f01  g1476 ( .o(n6964), .a(net_9935) );
in01f01  g1477 ( .o(n6965), .a(n6582) );
in01f01  g1478 ( .o(n6966_1), .a(n6606) );
oa22f01  g1479 ( .o(n6967), .a(n6966_1), .b(n6964), .c(n6965), .d(n6963) );
no04f01  g1480 ( .o(n6968), .a(n6967), .b(n6962_1), .c(n6960), .d(n6956) );
na04f01  g1481 ( .o(n755), .a(n6968), .b(n6953), .c(n6952), .d(n6951) );
in01f01  g1482 ( .o(n6970), .a(net_9748) );
no02f01  g1483 ( .o(n6971_1), .a(n5686), .b(n5672) );
in01f01  g1484 ( .o(n6972), .a(net_9739) );
in01f01  g1485 ( .o(n6973), .a(_net_9117) );
no02f01  g1486 ( .o(n6974), .a(n6973), .b(n6972) );
na03f01  g1487 ( .o(n6975), .a(n6971_1), .b(x4520), .c(x6599) );
no02f01  g1488 ( .o(n6976_1), .a(n6974), .b(n6971_1) );
na02f01  g1489 ( .o(n6977), .a(n6976_1), .b(x6599) );
oa12f01  g1490 ( .o(n760), .a(n6975), .b(n6977), .c(n6970) );
in01f01  g1491 ( .o(n6979), .a(x3828) );
in01f01  g1492 ( .o(n6980), .a(_net_10138) );
na02f01  g1493 ( .o(n6981_1), .a(n6980), .b(_net_10139) );
ao12f01  g1494 ( .o(n765), .a(n5658), .b(n6981_1), .c(n6979) );
in01f01  g1495 ( .o(n6983), .a(net_10514) );
no02f01  g1496 ( .o(n778), .a(n6164_1), .b(n6983) );
in01f01  g1497 ( .o(n6985_1), .a(net_10088) );
no04f01  g1498 ( .o(n6986), .a(n6559), .b(n5771), .c(n5664), .d(x6496) );
in01f01  g1499 ( .o(n6987), .a(n6986) );
na02f01  g1500 ( .o(n6988), .a(n6987), .b(x6599) );
na02f01  g1501 ( .o(n6989_1), .a(n6986), .b(x6599) );
oa22f01  g1502 ( .o(n783), .a(n6989_1), .b(n5516), .c(n6988), .d(n6985_1) );
in01f01  g1503 ( .o(n6991), .a(_net_10216) );
ao12f01  g1504 ( .o(n6992), .a(n5658), .b(n6887), .c(x5077) );
oa12f01  g1505 ( .o(n788), .a(n6992), .b(n6885_1), .c(n6991) );
in01f01  g1506 ( .o(n6994), .a(_net_10333) );
no02f01  g1507 ( .o(n6995), .a(n6994), .b(_net_10371) );
in01f01  g1508 ( .o(n6996), .a(_net_10371) );
no02f01  g1509 ( .o(n6997), .a(_net_10333), .b(n6996) );
in01f01  g1510 ( .o(n6998_1), .a(n6997) );
in01f01  g1511 ( .o(n6999), .a(_net_10332) );
no02f01  g1512 ( .o(n7000), .a(n6999), .b(_net_10370) );
ao12f01  g1513 ( .o(n7001), .a(n6995), .b(n7000), .c(n6998_1) );
in01f01  g1514 ( .o(n7002), .a(n7001) );
in01f01  g1515 ( .o(n7003_1), .a(_net_10370) );
no02f01  g1516 ( .o(n7004), .a(_net_10332), .b(n7003_1) );
in01f01  g1517 ( .o(n7005), .a(_net_10369) );
no02f01  g1518 ( .o(n7006), .a(n7005), .b(_net_10331) );
in01f01  g1519 ( .o(n7007_1), .a(_net_10368) );
no02f01  g1520 ( .o(n7008), .a(_net_10330), .b(n7007_1) );
in01f01  g1521 ( .o(n7009), .a(n7008) );
in01f01  g1522 ( .o(n7010), .a(_net_10367) );
no02f01  g1523 ( .o(n7011), .a(_net_10329), .b(n7010) );
in01f01  g1524 ( .o(n7012_1), .a(_net_10366) );
no02f01  g1525 ( .o(n7013), .a(_net_10328), .b(n7012_1) );
in01f01  g1526 ( .o(n7014), .a(n7013) );
in01f01  g1527 ( .o(n7015), .a(_net_10365) );
no02f01  g1528 ( .o(n7016), .a(n7015), .b(_net_10327) );
in01f01  g1529 ( .o(n7017_1), .a(_net_10327) );
in01f01  g1530 ( .o(n7018), .a(_net_10326) );
no02f01  g1531 ( .o(n7019), .a(_net_10364), .b(n7018) );
in01f01  g1532 ( .o(n7020), .a(n7019) );
oa12f01  g1533 ( .o(n7021_1), .a(n7017_1), .b(n7020), .c(_net_10365) );
oa12f01  g1534 ( .o(n7022), .a(_net_10365), .b(n7020), .c(n7017_1) );
na02f01  g1535 ( .o(n7023), .a(n7022), .b(n7021_1) );
in01f01  g1536 ( .o(n7024), .a(_net_10364) );
no02f01  g1537 ( .o(n7025), .a(n7024), .b(_net_10326) );
in01f01  g1538 ( .o(n7026_1), .a(n7025) );
in01f01  g1539 ( .o(n7027), .a(_net_10325) );
no02f01  g1540 ( .o(n7028), .a(n7027), .b(_net_10363) );
in01f01  g1541 ( .o(n7029), .a(_net_10362) );
no02f01  g1542 ( .o(n7030_1), .a(_net_10324), .b(n7029) );
in01f01  g1543 ( .o(n7031), .a(_net_10363) );
no02f01  g1544 ( .o(n7032), .a(_net_10325), .b(n7031) );
no02f01  g1545 ( .o(n7033), .a(n7032), .b(n7030_1) );
no02f01  g1546 ( .o(n7034_1), .a(n7033), .b(n7028) );
in01f01  g1547 ( .o(n7035), .a(n7034_1) );
na02f01  g1548 ( .o(n7036), .a(n7035), .b(n7026_1) );
oa12f01  g1549 ( .o(n7037), .a(n7023), .b(n7036), .c(n7016) );
na02f01  g1550 ( .o(n7038), .a(n7037), .b(n7014) );
no02f01  g1551 ( .o(n7039_1), .a(n7038), .b(n7011) );
na02f01  g1552 ( .o(n7040), .a(n7039_1), .b(n7009) );
in01f01  g1553 ( .o(n7041), .a(n7011) );
in01f01  g1554 ( .o(n7042), .a(_net_10329) );
no02f01  g1555 ( .o(n7043), .a(n7042), .b(_net_10367) );
in01f01  g1556 ( .o(n7044_1), .a(_net_10328) );
no02f01  g1557 ( .o(n7045), .a(n7044_1), .b(_net_10366) );
ao12f01  g1558 ( .o(n7046), .a(n7043), .b(n7045), .c(n7041) );
no02f01  g1559 ( .o(n7047), .a(n7046), .b(n7008) );
in01f01  g1560 ( .o(n7048_1), .a(_net_10331) );
in01f01  g1561 ( .o(n7049), .a(_net_10330) );
no02f01  g1562 ( .o(n7050), .a(n7049), .b(_net_10368) );
no02f01  g1563 ( .o(n7051), .a(_net_10369), .b(n7048_1) );
no02f01  g1564 ( .o(n7052), .a(n7051), .b(n7050) );
ao12f01  g1565 ( .o(n7053_1), .a(n7052), .b(n7006), .c(n7048_1) );
no02f01  g1566 ( .o(n7054), .a(n7053_1), .b(n7047) );
ao12f01  g1567 ( .o(n7055), .a(n7006), .b(n7054), .c(n7040) );
na02f01  g1568 ( .o(n7056), .a(n7053_1), .b(n7005) );
in01f01  g1569 ( .o(n7057), .a(n7056) );
no02f01  g1570 ( .o(n7058_1), .a(n7057), .b(n7055) );
no02f01  g1571 ( .o(n7059), .a(n7058_1), .b(n7004) );
na02f01  g1572 ( .o(n7060), .a(n7059), .b(n6998_1) );
in01f01  g1573 ( .o(n7061), .a(n7060) );
in01f01  g1574 ( .o(n7062), .a(_net_10372) );
no02f01  g1575 ( .o(n7063_1), .a(_net_10334), .b(n7062) );
in01f01  g1576 ( .o(n7064), .a(_net_10334) );
no02f01  g1577 ( .o(n7065), .a(n7064), .b(_net_10372) );
no02f01  g1578 ( .o(n7066), .a(n7065), .b(n7063_1) );
in01f01  g1579 ( .o(n7067), .a(n7066) );
oa12f01  g1580 ( .o(n7068_1), .a(n7067), .b(n7061), .c(n7002) );
na03f01  g1581 ( .o(n7069), .a(n7066), .b(n7060), .c(n7001) );
na02f01  g1582 ( .o(n793), .a(n7069), .b(n7068_1) );
in01f01  g1583 ( .o(n7071), .a(_net_170) );
in01f01  g1584 ( .o(n7072), .a(n5941) );
in01f01  g1585 ( .o(n7073_1), .a(_net_9293) );
no02f01  g1586 ( .o(n7074), .a(n6026), .b(n7073_1) );
ao12f01  g1587 ( .o(n7075), .a(n7074), .b(n6028_1), .c(n7072) );
oa12f01  g1588 ( .o(n798), .a(n7075), .b(n6022), .c(n7071) );
in01f01  g1589 ( .o(n7077), .a(_net_10205) );
ao12f01  g1590 ( .o(n7078_1), .a(n5658), .b(n6887), .c(x5790) );
oa12f01  g1591 ( .o(n803), .a(n7078_1), .b(n6885_1), .c(n7077) );
na02f01  g1592 ( .o(n7080), .a(n6056), .b(net_258) );
na02f01  g1593 ( .o(n7081), .a(n6055), .b(net_9986) );
ao22f01  g1594 ( .o(n7082_1), .a(n6062_1), .b(x4209), .c(n6060), .d(_net_10437) );
na04f01  g1595 ( .o(n808), .a(n7082_1), .b(n7081), .c(n7080), .d(n6058) );
ao12f01  g1596 ( .o(n7084), .a(n5658), .b(n6875_1), .c(net_236) );
ao22f01  g1597 ( .o(n7085), .a(n6878), .b(x5790), .c(n6877), .d(net_9897) );
na02f01  g1598 ( .o(n813), .a(n7085), .b(n7084) );
no02f01  g1599 ( .o(n7087), .a(_net_9376), .b(_net_9375) );
in01f01  g1600 ( .o(n7088), .a(_net_9375) );
in01f01  g1601 ( .o(n7089), .a(_net_9376) );
no02f01  g1602 ( .o(n7090), .a(n7089), .b(n7088) );
no02f01  g1603 ( .o(n7091_1), .a(n7090), .b(n7087) );
no02f01  g1604 ( .o(n7092), .a(n7091_1), .b(_net_9377) );
in01f01  g1605 ( .o(n7093), .a(n7091_1) );
no02f01  g1606 ( .o(n7094), .a(n7093), .b(n6106) );
in01f01  g1607 ( .o(n7095_1), .a(_net_9371) );
no02f01  g1608 ( .o(n7096), .a(_net_9372), .b(n7095_1) );
in01f01  g1609 ( .o(n7097), .a(_net_9372) );
no02f01  g1610 ( .o(n7098), .a(n7097), .b(_net_9371) );
no02f01  g1611 ( .o(n7099), .a(n7098), .b(n7096) );
in01f01  g1612 ( .o(n7100_1), .a(n7099) );
no03f01  g1613 ( .o(n7101), .a(n7100_1), .b(n7094), .c(n7092) );
no02f01  g1614 ( .o(n7102), .a(n7094), .b(n7092) );
no02f01  g1615 ( .o(n7103), .a(n7099), .b(n7102) );
in01f01  g1616 ( .o(n7104_1), .a(_net_9374) );
no02f01  g1617 ( .o(n7105), .a(_net_9373), .b(n7104_1) );
in01f01  g1618 ( .o(n7106), .a(_net_9373) );
no02f01  g1619 ( .o(n7107), .a(n7106), .b(_net_9374) );
no02f01  g1620 ( .o(n7108_1), .a(n7107), .b(n7105) );
no02f01  g1621 ( .o(n7109), .a(n7108_1), .b(_net_9370) );
in01f01  g1622 ( .o(n7110), .a(_net_9370) );
in01f01  g1623 ( .o(n7111), .a(n7108_1) );
no02f01  g1624 ( .o(n7112), .a(n7111), .b(n7110) );
no02f01  g1625 ( .o(n7113_1), .a(n7112), .b(n7109) );
in01f01  g1626 ( .o(n7114), .a(n7113_1) );
no03f01  g1627 ( .o(n7115), .a(n7114), .b(n7103), .c(n7101) );
no02f01  g1628 ( .o(n7116), .a(n7103), .b(n7101) );
no02f01  g1629 ( .o(n7117), .a(n7113_1), .b(n7116) );
no02f01  g1630 ( .o(n7118_1), .a(n7117), .b(n7115) );
in01f01  g1631 ( .o(n7119), .a(net_9493) );
na02f01  g1632 ( .o(n7120), .a(n6081), .b(n6075) );
no03f01  g1633 ( .o(n7121), .a(n7120), .b(n6089), .c(n7119) );
in01f01  g1634 ( .o(n7122), .a(net_9501) );
na02f01  g1635 ( .o(n7123_1), .a(n6081), .b(n6084) );
no03f01  g1636 ( .o(n7124), .a(n7123_1), .b(n6089), .c(n7122) );
no02f01  g1637 ( .o(n7125), .a(n7120), .b(n6071) );
na02f01  g1638 ( .o(n7126), .a(n7125), .b(net_9477) );
no02f01  g1639 ( .o(n7127), .a(n7123_1), .b(n6071) );
na02f01  g1640 ( .o(n7128_1), .a(n7127), .b(net_9485) );
na02f01  g1641 ( .o(n7129), .a(n7128_1), .b(n7126) );
na02f01  g1642 ( .o(n7130), .a(n6097), .b(n6075) );
no02f01  g1643 ( .o(n7131), .a(n7130), .b(n6071) );
na02f01  g1644 ( .o(n7132), .a(n6097), .b(n6084) );
no02f01  g1645 ( .o(n7133_1), .a(n7132), .b(n6071) );
ao22f01  g1646 ( .o(n7134), .a(n7133_1), .b(net_9453), .c(n7131), .d(net_9445) );
no02f01  g1647 ( .o(n7135), .a(n7130), .b(n6089) );
no02f01  g1648 ( .o(n7136), .a(n7132), .b(n6089) );
ao22f01  g1649 ( .o(n7137), .a(n7136), .b(net_9469), .c(n7135), .d(net_9461) );
na02f01  g1650 ( .o(n7138_1), .a(n7137), .b(n7134) );
no04f01  g1651 ( .o(n7139), .a(n7138_1), .b(n7129), .c(n7124), .d(n7121) );
in01f01  g1652 ( .o(n7140), .a(n7139) );
na04f01  g1653 ( .o(n7141), .a(n6097), .b(n6075), .c(n6089), .d(net_9439) );
na04f01  g1654 ( .o(n7142), .a(n6097), .b(n6084), .c(n6089), .d(net_9447) );
na04f01  g1655 ( .o(n7143_1), .a(n6097), .b(n6075), .c(n6071), .d(net_9455) );
na04f01  g1656 ( .o(n7144), .a(n6097), .b(n6084), .c(n6071), .d(net_9463) );
na04f01  g1657 ( .o(n7145), .a(n7144), .b(n7143_1), .c(n7142), .d(n7141) );
na04f01  g1658 ( .o(n7146), .a(n6081), .b(n6084), .c(n6071), .d(net_9495) );
na04f01  g1659 ( .o(n7147), .a(n6081), .b(n6075), .c(n6071), .d(net_9487) );
na04f01  g1660 ( .o(n7148_1), .a(n6081), .b(n6084), .c(n6089), .d(net_9479) );
na04f01  g1661 ( .o(n7149), .a(n6081), .b(n6075), .c(n6089), .d(net_9471) );
na04f01  g1662 ( .o(n7150), .a(n7149), .b(n7148_1), .c(n7147), .d(n7146) );
no02f01  g1663 ( .o(n7151), .a(n7150), .b(n7145) );
na02f01  g1664 ( .o(n7152), .a(n7151), .b(n6128) );
in01f01  g1665 ( .o(n7153_1), .a(net_9439) );
no04f01  g1666 ( .o(n7154), .a(n6081), .b(n6084), .c(n6071), .d(n7153_1) );
in01f01  g1667 ( .o(n7155), .a(net_9447) );
no04f01  g1668 ( .o(n7156), .a(n6081), .b(n6075), .c(n6071), .d(n7155) );
in01f01  g1669 ( .o(n7157), .a(net_9455) );
no04f01  g1670 ( .o(n7158_1), .a(n6081), .b(n6084), .c(n6089), .d(n7157) );
in01f01  g1671 ( .o(n7159), .a(net_9463) );
no04f01  g1672 ( .o(n7160), .a(n6081), .b(n6075), .c(n6089), .d(n7159) );
no04f01  g1673 ( .o(n7161), .a(n7160), .b(n7158_1), .c(n7156), .d(n7154) );
in01f01  g1674 ( .o(n7162), .a(net_9495) );
no04f01  g1675 ( .o(n7163_1), .a(n6097), .b(n6075), .c(n6089), .d(n7162) );
in01f01  g1676 ( .o(n7164), .a(net_9487) );
no04f01  g1677 ( .o(n7165), .a(n6097), .b(n6084), .c(n6089), .d(n7164) );
in01f01  g1678 ( .o(n7166), .a(net_9479) );
no04f01  g1679 ( .o(n7167), .a(n6097), .b(n6075), .c(n6071), .d(n7166) );
in01f01  g1680 ( .o(n7168_1), .a(net_9471) );
no04f01  g1681 ( .o(n7169), .a(n6097), .b(n6084), .c(n6071), .d(n7168_1) );
no04f01  g1682 ( .o(n7170), .a(n7169), .b(n7167), .c(n7165), .d(n7163_1) );
na02f01  g1683 ( .o(n7171), .a(n7170), .b(n7161) );
na02f01  g1684 ( .o(n7172), .a(n7171), .b(n6103) );
na02f01  g1685 ( .o(n7173_1), .a(n7172), .b(n7152) );
in01f01  g1686 ( .o(n7174), .a(net_9444) );
no04f01  g1687 ( .o(n7175), .a(n6081), .b(n6084), .c(n6071), .d(n7174) );
in01f01  g1688 ( .o(n7176), .a(net_9452) );
no04f01  g1689 ( .o(n7177_1), .a(n6081), .b(n6075), .c(n6071), .d(n7176) );
in01f01  g1690 ( .o(n7178), .a(net_9500) );
no04f01  g1691 ( .o(n7179), .a(n6097), .b(n6075), .c(n6089), .d(n7178) );
in01f01  g1692 ( .o(n7180), .a(net_9492) );
no04f01  g1693 ( .o(n7181), .a(n6097), .b(n6084), .c(n6089), .d(n7180) );
no04f01  g1694 ( .o(n7182_1), .a(n7181), .b(n7179), .c(n7177_1), .d(n7175) );
in01f01  g1695 ( .o(n7183), .a(net_9484) );
no04f01  g1696 ( .o(n7184), .a(n6097), .b(n6075), .c(n6071), .d(n7183) );
in01f01  g1697 ( .o(n7185), .a(net_9476) );
no04f01  g1698 ( .o(n7186), .a(n6097), .b(n6084), .c(n6071), .d(n7185) );
in01f01  g1699 ( .o(n7187_1), .a(net_9460) );
no04f01  g1700 ( .o(n7188), .a(n6081), .b(n6084), .c(n6089), .d(n7187_1) );
in01f01  g1701 ( .o(n7189), .a(net_9468) );
no04f01  g1702 ( .o(n7190), .a(n6081), .b(n6075), .c(n6089), .d(n7189) );
no04f01  g1703 ( .o(n7191), .a(n7190), .b(n7188), .c(n7186), .d(n7184) );
na02f01  g1704 ( .o(n7192_1), .a(n7191), .b(n7182_1) );
na04f01  g1705 ( .o(n7193), .a(n6081), .b(n6075), .c(n6089), .d(net_9475) );
na04f01  g1706 ( .o(n7194), .a(n6081), .b(n6084), .c(n6089), .d(net_9483) );
na04f01  g1707 ( .o(n7195), .a(n6081), .b(n6084), .c(n6071), .d(net_9499) );
na04f01  g1708 ( .o(n7196), .a(n6081), .b(n6075), .c(n6071), .d(net_9491) );
na04f01  g1709 ( .o(n7197_1), .a(n7196), .b(n7195), .c(n7194), .d(n7193) );
na04f01  g1710 ( .o(n7198), .a(n6097), .b(n6084), .c(n6071), .d(net_9467) );
na04f01  g1711 ( .o(n7199), .a(n6097), .b(n6075), .c(n6071), .d(net_9459) );
na04f01  g1712 ( .o(n7200), .a(n6097), .b(n6075), .c(n6089), .d(net_9443) );
na04f01  g1713 ( .o(n7201), .a(n6097), .b(n6084), .c(n6089), .d(net_9451) );
na04f01  g1714 ( .o(n7202_1), .a(n7201), .b(n7200), .c(n7199), .d(n7198) );
no02f01  g1715 ( .o(n7203), .a(n7202_1), .b(n7197_1) );
no02f01  g1716 ( .o(n7204), .a(n7203), .b(n7192_1) );
na04f01  g1717 ( .o(n7205), .a(n6097), .b(n6075), .c(n6089), .d(net_9444) );
na04f01  g1718 ( .o(n7206_1), .a(n6097), .b(n6084), .c(n6089), .d(net_9452) );
na04f01  g1719 ( .o(n7207), .a(n6081), .b(n6084), .c(n6071), .d(net_9500) );
na04f01  g1720 ( .o(n7208), .a(n6081), .b(n6075), .c(n6071), .d(net_9492) );
na04f01  g1721 ( .o(n7209), .a(n7208), .b(n7207), .c(n7206_1), .d(n7205) );
na04f01  g1722 ( .o(n7210), .a(n6081), .b(n6084), .c(n6089), .d(net_9484) );
na04f01  g1723 ( .o(n7211_1), .a(n6081), .b(n6075), .c(n6089), .d(net_9476) );
na04f01  g1724 ( .o(n7212), .a(n6097), .b(n6075), .c(n6071), .d(net_9460) );
na04f01  g1725 ( .o(n7213), .a(n6097), .b(n6084), .c(n6071), .d(net_9468) );
na04f01  g1726 ( .o(n7214), .a(n7213), .b(n7212), .c(n7211_1), .d(n7210) );
no02f01  g1727 ( .o(n7215), .a(n7214), .b(n7209) );
in01f01  g1728 ( .o(n7216_1), .a(net_9475) );
no04f01  g1729 ( .o(n7217), .a(n6097), .b(n6084), .c(n6071), .d(n7216_1) );
in01f01  g1730 ( .o(n7218), .a(net_9483) );
no04f01  g1731 ( .o(n7219), .a(n6097), .b(n6075), .c(n6071), .d(n7218) );
in01f01  g1732 ( .o(n7220), .a(net_9499) );
no04f01  g1733 ( .o(n7221_1), .a(n6097), .b(n6075), .c(n6089), .d(n7220) );
in01f01  g1734 ( .o(n7222), .a(net_9491) );
no04f01  g1735 ( .o(n7223), .a(n6097), .b(n6084), .c(n6089), .d(n7222) );
no04f01  g1736 ( .o(n7224), .a(n7223), .b(n7221_1), .c(n7219), .d(n7217) );
in01f01  g1737 ( .o(n7225), .a(net_9467) );
no04f01  g1738 ( .o(n7226_1), .a(n6081), .b(n6075), .c(n6089), .d(n7225) );
in01f01  g1739 ( .o(n7227), .a(net_9459) );
no04f01  g1740 ( .o(n7228), .a(n6081), .b(n6084), .c(n6089), .d(n7227) );
in01f01  g1741 ( .o(n7229), .a(net_9443) );
no04f01  g1742 ( .o(n7230), .a(n6081), .b(n6084), .c(n6071), .d(n7229) );
in01f01  g1743 ( .o(n7231_1), .a(net_9451) );
no04f01  g1744 ( .o(n7232), .a(n6081), .b(n6075), .c(n6071), .d(n7231_1) );
no04f01  g1745 ( .o(n7233), .a(n7232), .b(n7230), .c(n7228), .d(n7226_1) );
na02f01  g1746 ( .o(n7234), .a(n7233), .b(n7224) );
no02f01  g1747 ( .o(n7235_1), .a(n7234), .b(n7215) );
no02f01  g1748 ( .o(n7236), .a(n7235_1), .b(n7204) );
no02f01  g1749 ( .o(n7237), .a(n7236), .b(n7173_1) );
no02f01  g1750 ( .o(n7238), .a(n7171), .b(n6103) );
no02f01  g1751 ( .o(n7239), .a(n7151), .b(n6128) );
no02f01  g1752 ( .o(n7240_1), .a(n7239), .b(n7238) );
na02f01  g1753 ( .o(n7241), .a(n7234), .b(n7215) );
na02f01  g1754 ( .o(n7242), .a(n7203), .b(n7192_1) );
na02f01  g1755 ( .o(n7243), .a(n7242), .b(n7241) );
no02f01  g1756 ( .o(n7244), .a(n7243), .b(n7240_1) );
in01f01  g1757 ( .o(n7245_1), .a(net_9465) );
no04f01  g1758 ( .o(n7246), .a(n6081), .b(n6075), .c(n6089), .d(n7245_1) );
in01f01  g1759 ( .o(n7247), .a(net_9457) );
no04f01  g1760 ( .o(n7248), .a(n6081), .b(n6084), .c(n6089), .d(n7247) );
in01f01  g1761 ( .o(n7249), .a(net_9441) );
no04f01  g1762 ( .o(n7250_1), .a(n6081), .b(n6084), .c(n6071), .d(n7249) );
in01f01  g1763 ( .o(n7251), .a(net_9449) );
no04f01  g1764 ( .o(n7252), .a(n6081), .b(n6075), .c(n6071), .d(n7251) );
no04f01  g1765 ( .o(n7253), .a(n7252), .b(n7250_1), .c(n7248), .d(n7246) );
in01f01  g1766 ( .o(n7254), .a(net_9497) );
no04f01  g1767 ( .o(n7255_1), .a(n6097), .b(n6075), .c(n6089), .d(n7254) );
in01f01  g1768 ( .o(n7256), .a(net_9489) );
no04f01  g1769 ( .o(n7257), .a(n6097), .b(n6084), .c(n6089), .d(n7256) );
in01f01  g1770 ( .o(n7258), .a(net_9481) );
no04f01  g1771 ( .o(n7259), .a(n6097), .b(n6075), .c(n6071), .d(n7258) );
in01f01  g1772 ( .o(n7260_1), .a(net_9473) );
no04f01  g1773 ( .o(n7261), .a(n6097), .b(n6084), .c(n6071), .d(n7260_1) );
no04f01  g1774 ( .o(n7262), .a(n7261), .b(n7259), .c(n7257), .d(n7255_1) );
na02f01  g1775 ( .o(n7263), .a(n7262), .b(n7253) );
na04f01  g1776 ( .o(n7264), .a(n6081), .b(n6084), .c(n6071), .d(net_9498) );
na04f01  g1777 ( .o(n7265_1), .a(n6081), .b(n6075), .c(n6071), .d(net_9490) );
na04f01  g1778 ( .o(n7266), .a(n6081), .b(n6084), .c(n6089), .d(net_9482) );
na04f01  g1779 ( .o(n7267), .a(n6081), .b(n6075), .c(n6089), .d(net_9474) );
na04f01  g1780 ( .o(n7268), .a(n7267), .b(n7266), .c(n7265_1), .d(n7264) );
na04f01  g1781 ( .o(n7269), .a(n6097), .b(n6075), .c(n6089), .d(net_9442) );
na04f01  g1782 ( .o(n7270_1), .a(n6097), .b(n6084), .c(n6089), .d(net_9450) );
na04f01  g1783 ( .o(n7271), .a(n6097), .b(n6084), .c(n6071), .d(net_9466) );
na04f01  g1784 ( .o(n7272), .a(n6097), .b(n6075), .c(n6071), .d(net_9458) );
na04f01  g1785 ( .o(n7273), .a(n7272), .b(n7271), .c(n7270_1), .d(n7269) );
no02f01  g1786 ( .o(n7274), .a(n7273), .b(n7268) );
no02f01  g1787 ( .o(n7275_1), .a(n7274), .b(n7263) );
na04f01  g1788 ( .o(n7276), .a(n6097), .b(n6084), .c(n6071), .d(net_9465) );
na04f01  g1789 ( .o(n7277), .a(n6097), .b(n6075), .c(n6071), .d(net_9457) );
na04f01  g1790 ( .o(n7278), .a(n6097), .b(n6075), .c(n6089), .d(net_9441) );
na04f01  g1791 ( .o(n7279), .a(n6097), .b(n6084), .c(n6089), .d(net_9449) );
na04f01  g1792 ( .o(n7280_1), .a(n7279), .b(n7278), .c(n7277), .d(n7276) );
na04f01  g1793 ( .o(n7281), .a(n6081), .b(n6084), .c(n6071), .d(net_9497) );
na04f01  g1794 ( .o(n7282), .a(n6081), .b(n6075), .c(n6071), .d(net_9489) );
na04f01  g1795 ( .o(n7283), .a(n6081), .b(n6084), .c(n6089), .d(net_9481) );
na04f01  g1796 ( .o(n7284), .a(n6081), .b(n6075), .c(n6089), .d(net_9473) );
na04f01  g1797 ( .o(n7285_1), .a(n7284), .b(n7283), .c(n7282), .d(n7281) );
no02f01  g1798 ( .o(n7286), .a(n7285_1), .b(n7280_1) );
in01f01  g1799 ( .o(n7287), .a(net_9498) );
no04f01  g1800 ( .o(n7288), .a(n6097), .b(n6075), .c(n6089), .d(n7287) );
in01f01  g1801 ( .o(n7289), .a(net_9490) );
no04f01  g1802 ( .o(n7290_1), .a(n6097), .b(n6084), .c(n6089), .d(n7289) );
in01f01  g1803 ( .o(n7291), .a(net_9482) );
no04f01  g1804 ( .o(n7292), .a(n6097), .b(n6075), .c(n6071), .d(n7291) );
in01f01  g1805 ( .o(n7293), .a(net_9474) );
no04f01  g1806 ( .o(n7294), .a(n6097), .b(n6084), .c(n6071), .d(n7293) );
no04f01  g1807 ( .o(n7295_1), .a(n7294), .b(n7292), .c(n7290_1), .d(n7288) );
in01f01  g1808 ( .o(n7296), .a(net_9442) );
no04f01  g1809 ( .o(n7297), .a(n6081), .b(n6084), .c(n6071), .d(n7296) );
in01f01  g1810 ( .o(n7298), .a(net_9450) );
no04f01  g1811 ( .o(n7299), .a(n6081), .b(n6075), .c(n6071), .d(n7298) );
in01f01  g1812 ( .o(n7300_1), .a(net_9466) );
no04f01  g1813 ( .o(n7301), .a(n6081), .b(n6075), .c(n6089), .d(n7300_1) );
in01f01  g1814 ( .o(n7302), .a(net_9458) );
no04f01  g1815 ( .o(n7303), .a(n6081), .b(n6084), .c(n6089), .d(n7302) );
no04f01  g1816 ( .o(n7304_1), .a(n7303), .b(n7301), .c(n7299), .d(n7297) );
na02f01  g1817 ( .o(n7305), .a(n7304_1), .b(n7295_1) );
no02f01  g1818 ( .o(n7306), .a(n7305), .b(n7286) );
no02f01  g1819 ( .o(n7307), .a(n7120), .b(n6089) );
no02f01  g1820 ( .o(n7308_1), .a(n7123_1), .b(n6089) );
ao22f01  g1821 ( .o(n7309), .a(n7308_1), .b(net_9496), .c(n7307), .d(net_9488) );
ao22f01  g1822 ( .o(n7310), .a(n7127), .b(net_9480), .c(n7125), .d(net_9472) );
na02f01  g1823 ( .o(n7311), .a(n7310), .b(n7309) );
ao22f01  g1824 ( .o(n7312_1), .a(n7133_1), .b(net_9448), .c(n7131), .d(net_9440) );
ao22f01  g1825 ( .o(n7313), .a(n7136), .b(net_9464), .c(n7135), .d(net_9456) );
na02f01  g1826 ( .o(n7314), .a(n7313), .b(n7312_1) );
no02f01  g1827 ( .o(n7315), .a(n7314), .b(n7311) );
no03f01  g1828 ( .o(n7316), .a(n7315), .b(n7306), .c(n7275_1) );
na02f01  g1829 ( .o(n7317_1), .a(n7305), .b(n7286) );
na02f01  g1830 ( .o(n7318), .a(n7274), .b(n7263) );
na04f01  g1831 ( .o(n7319), .a(n7313), .b(n7312_1), .c(n7310), .d(n7309) );
ao12f01  g1832 ( .o(n7320), .a(n7319), .b(n7318), .c(n7317_1) );
no02f01  g1833 ( .o(n7321_1), .a(n7320), .b(n7316) );
no03f01  g1834 ( .o(n7322), .a(n7321_1), .b(n7244), .c(n7237) );
na02f01  g1835 ( .o(n7323), .a(n7243), .b(n7240_1) );
na02f01  g1836 ( .o(n7324), .a(n7236), .b(n7173_1) );
na03f01  g1837 ( .o(n7325), .a(n7319), .b(n7318), .c(n7317_1) );
oa12f01  g1838 ( .o(n7326_1), .a(n7315), .b(n7306), .c(n7275_1) );
na02f01  g1839 ( .o(n7327), .a(n7326_1), .b(n7325) );
ao12f01  g1840 ( .o(n7328), .a(n7327), .b(n7324), .c(n7323) );
no02f01  g1841 ( .o(n7329), .a(n7328), .b(n7322) );
no02f01  g1842 ( .o(n7330), .a(n7329), .b(n7140) );
na03f01  g1843 ( .o(n7331_1), .a(n7327), .b(n7324), .c(n7323) );
oa12f01  g1844 ( .o(n7332), .a(n7321_1), .b(n7244), .c(n7237) );
na02f01  g1845 ( .o(n7333), .a(n7332), .b(n7331_1) );
no02f01  g1846 ( .o(n7334), .a(n7333), .b(n7139) );
no02f01  g1847 ( .o(n7335), .a(n7334), .b(n7330) );
no02f01  g1848 ( .o(n7336_1), .a(n7335), .b(n7118_1) );
in01f01  g1849 ( .o(n7337), .a(n7118_1) );
na02f01  g1850 ( .o(n7338), .a(n7333), .b(n7139) );
na02f01  g1851 ( .o(n7339), .a(n7329), .b(n7140) );
na02f01  g1852 ( .o(n7340), .a(n7339), .b(n7338) );
no02f01  g1853 ( .o(n7341_1), .a(n7340), .b(n7337) );
oa12f01  g1854 ( .o(n7342), .a(n6148), .b(n7341_1), .c(n7336_1) );
ao12f01  g1855 ( .o(n7343), .a(n6131_1), .b(n6147), .c(_net_9362) );
na02f01  g1856 ( .o(n818), .a(n7343), .b(n7342) );
in01f01  g1857 ( .o(n7345), .a(n6160_1) );
no02f01  g1858 ( .o(n7346_1), .a(n6743_1), .b(n6159) );
in01f01  g1859 ( .o(n7347), .a(n7346_1) );
in01f01  g1860 ( .o(n7348), .a(n6159) );
na04f01  g1861 ( .o(n7349), .a(n7348), .b(_net_133), .c(n6031), .d(net_10175) );
no02f01  g1862 ( .o(n7350), .a(n6160_1), .b(n5658) );
na03f01  g1863 ( .o(n7351_1), .a(n7350), .b(n7349), .c(n7347) );
in01f01  g1864 ( .o(n7352), .a(n7351_1) );
no02f01  g1865 ( .o(n7353), .a(n7352), .b(n7345) );
na02f01  g1866 ( .o(n7354), .a(n7353), .b(x5647) );
na02f01  g1867 ( .o(n7355_1), .a(n7351_1), .b(n5658) );
na02f01  g1868 ( .o(n7356), .a(n7352), .b(net_9669) );
no02f01  g1869 ( .o(n7357), .a(n7352), .b(n7347) );
no02f01  g1870 ( .o(n7358), .a(n7352), .b(n7349) );
ao22f01  g1871 ( .o(n7359), .a(n7358), .b(net_238), .c(n7357), .d(_net_10102) );
na04f01  g1872 ( .o(n823), .a(n7359), .b(n7356), .c(n7355_1), .d(n7354) );
in01f01  g1873 ( .o(n7361), .a(_net_10431) );
ao12f01  g1874 ( .o(n7362), .a(n5658), .b(n6052_1), .c(x4694) );
oa12f01  g1875 ( .o(n828), .a(n7362), .b(n6048), .c(n7361) );
in01f01  g1876 ( .o(n7364), .a(net_9749) );
na02f01  g1877 ( .o(n7365_1), .a(n6971_1), .b(x6599) );
in01f01  g1878 ( .o(n7366), .a(n6971_1) );
na02f01  g1879 ( .o(n7367), .a(n7366), .b(x6599) );
oa22f01  g1880 ( .o(n833), .a(n7367), .b(n7364), .c(n7365_1), .d(n5597_1) );
in01f01  g1881 ( .o(n7369), .a(_net_10478) );
in01f01  g1882 ( .o(n7370_1), .a(_net_10477) );
in01f01  g1883 ( .o(n7371), .a(_net_10476) );
in01f01  g1884 ( .o(n7372), .a(_net_10033) );
in01f01  g1885 ( .o(n7373), .a(_net_10475) );
no02f01  g1886 ( .o(n7374), .a(n7373), .b(n7372) );
no02f01  g1887 ( .o(n7375_1), .a(_net_10475), .b(_net_10033) );
in01f01  g1888 ( .o(n7376), .a(n7375_1) );
in01f01  g1889 ( .o(n7377), .a(_net_10474) );
no02f01  g1890 ( .o(n7378), .a(_net_10032), .b(_net_10474) );
in01f01  g1891 ( .o(n7379_1), .a(_net_10031) );
in01f01  g1892 ( .o(n7380), .a(_net_10473) );
no02f01  g1893 ( .o(n7381), .a(n7380), .b(n7379_1) );
in01f01  g1894 ( .o(n7382), .a(_net_10032) );
no02f01  g1895 ( .o(n7383), .a(n7382), .b(n7377) );
na02f01  g1896 ( .o(n7384_1), .a(n7382), .b(n7377) );
oa12f01  g1897 ( .o(n7385), .a(n7384_1), .b(n7383), .c(n7381) );
no02f01  g1898 ( .o(n7386), .a(_net_10028), .b(_net_10470) );
in01f01  g1899 ( .o(n7387), .a(n7386) );
in01f01  g1900 ( .o(n7388), .a(_net_10469) );
in01f01  g1901 ( .o(n7389_1), .a(_net_10027) );
no02f01  g1902 ( .o(n7390), .a(n7389_1), .b(n7388) );
ao12f01  g1903 ( .o(n7391), .a(_net_10470), .b(n7390), .c(_net_10028) );
ao12f01  g1904 ( .o(n7392), .a(_net_10028), .b(n7390), .c(_net_10470) );
no02f01  g1905 ( .o(n7393), .a(n7392), .b(n7391) );
no02f01  g1906 ( .o(n7394_1), .a(_net_10027), .b(_net_10469) );
in01f01  g1907 ( .o(n7395), .a(_net_10468) );
in01f01  g1908 ( .o(n7396), .a(_net_10026) );
no02f01  g1909 ( .o(n7397), .a(n7396), .b(n7395) );
in01f01  g1910 ( .o(n7398_1), .a(_net_10467) );
in01f01  g1911 ( .o(n7399), .a(_net_10025) );
no02f01  g1912 ( .o(n7400), .a(n7399), .b(n7398_1) );
no02f01  g1913 ( .o(n7401), .a(_net_10026), .b(_net_10468) );
in01f01  g1914 ( .o(n7402), .a(n7401) );
ao12f01  g1915 ( .o(n7403_1), .a(n7397), .b(n7402), .c(n7400) );
no02f01  g1916 ( .o(n7404), .a(n7403_1), .b(n7394_1) );
ao12f01  g1917 ( .o(n7405), .a(n7393), .b(n7404), .c(n7387) );
no02f01  g1918 ( .o(n7406), .a(_net_10471), .b(_net_10029) );
no02f01  g1919 ( .o(n7407), .a(_net_10473), .b(_net_10031) );
no02f01  g1920 ( .o(n7408_1), .a(_net_10472), .b(_net_10030) );
no04f01  g1921 ( .o(n7409), .a(n7408_1), .b(n7407), .c(n7406), .d(n7405) );
in01f01  g1922 ( .o(n7410), .a(n7407) );
in01f01  g1923 ( .o(n7411), .a(n7408_1) );
in01f01  g1924 ( .o(n7412), .a(_net_10030) );
in01f01  g1925 ( .o(n7413_1), .a(_net_10472) );
no02f01  g1926 ( .o(n7414), .a(n7413_1), .b(n7412) );
in01f01  g1927 ( .o(n7415), .a(_net_10471) );
no02f01  g1928 ( .o(n7416), .a(n7415), .b(n5897) );
ao12f01  g1929 ( .o(n7417), .a(n7414), .b(n7416), .c(n7411) );
in01f01  g1930 ( .o(n7418_1), .a(n7417) );
na02f01  g1931 ( .o(n7419), .a(n7418_1), .b(n7410) );
na02f01  g1932 ( .o(n7420), .a(n7385), .b(n7419) );
no02f01  g1933 ( .o(n7421), .a(n7420), .b(n7409) );
oa22f01  g1934 ( .o(n7422), .a(n7421), .b(n7378), .c(n7385), .d(n7377) );
ao12f01  g1935 ( .o(n7423_1), .a(n7374), .b(n7422), .c(n7376) );
no02f01  g1936 ( .o(n7424), .a(n7423_1), .b(n7371) );
in01f01  g1937 ( .o(n7425), .a(n7424) );
no02f01  g1938 ( .o(n7426), .a(n7425), .b(n7370_1) );
in01f01  g1939 ( .o(n7427), .a(n7426) );
no02f01  g1940 ( .o(n7428_1), .a(n7427), .b(n7369) );
in01f01  g1941 ( .o(n7429), .a(_net_10037) );
oa12f01  g1942 ( .o(n7430), .a(net_10490), .b(n6165), .c(_net_8831) );
no03f01  g1943 ( .o(n7431), .a(n7430), .b(n7429), .c(net_10514) );
oa12f01  g1944 ( .o(n7432_1), .a(n7431), .b(n7426), .c(_net_10478) );
in01f01  g1945 ( .o(n7433), .a(_net_10470) );
no02f01  g1946 ( .o(n7434), .a(_net_10468), .b(_net_10467) );
in01f01  g1947 ( .o(n7435), .a(n7434) );
no02f01  g1948 ( .o(n7436_1), .a(n7435), .b(_net_10469) );
na02f01  g1949 ( .o(n7437), .a(n7436_1), .b(n7433) );
no02f01  g1950 ( .o(n7438), .a(n7437), .b(_net_10471) );
in01f01  g1951 ( .o(n7439), .a(n7438) );
no02f01  g1952 ( .o(n7440), .a(n7439), .b(_net_10472) );
in01f01  g1953 ( .o(n7441_1), .a(n7440) );
no02f01  g1954 ( .o(n7442), .a(n7441_1), .b(_net_10473) );
in01f01  g1955 ( .o(n7443), .a(n7442) );
no02f01  g1956 ( .o(n7444), .a(n7443), .b(_net_10474) );
na02f01  g1957 ( .o(n7445), .a(n7444), .b(n7373) );
no02f01  g1958 ( .o(n7446_1), .a(n7445), .b(_net_10476) );
na03f01  g1959 ( .o(n7447), .a(n7446_1), .b(n7370_1), .c(_net_10478) );
ao12f01  g1960 ( .o(n7448), .a(_net_10478), .b(n7446_1), .c(n7370_1) );
in01f01  g1961 ( .o(n7449), .a(n7430) );
no02f01  g1962 ( .o(n7450), .a(n7429), .b(n6983) );
in01f01  g1963 ( .o(n7451_1), .a(n7450) );
no02f01  g1964 ( .o(n7452), .a(n7451_1), .b(n7448) );
no03f01  g1965 ( .o(n7453), .a(n7449), .b(n7429), .c(net_10514) );
ao22f01  g1966 ( .o(n7454), .a(n7453), .b(_net_10478), .c(n7452), .d(n7447) );
oa12f01  g1967 ( .o(n838), .a(n7454), .b(n7432_1), .c(n7428_1) );
ao12f01  g1968 ( .o(n7456), .a(n5658), .b(n5678), .c(_net_261) );
ao22f01  g1969 ( .o(n7457), .a(n5681_1), .b(x3949), .c(n5680), .d(net_9724) );
na02f01  g1970 ( .o(n843), .a(n7457), .b(n7456) );
ao22f01  g1971 ( .o(n7459), .a(n5842), .b(net_9749), .c(n5841), .d(_net_185) );
na02f01  g1972 ( .o(n7460_1), .a(n5847), .b(net_10046) );
ao22f01  g1973 ( .o(n7461), .a(n5850), .b(net_9848), .c(n5849_1), .d(net_9947) );
na03f01  g1974 ( .o(n848), .a(n7461), .b(n7460_1), .c(n7459) );
in01f01  g1975 ( .o(n7463), .a(net_10502) );
no02f01  g1976 ( .o(n7464), .a(n6570), .b(n5658) );
no02f01  g1977 ( .o(n7465_1), .a(n7464), .b(n6047_1) );
no02f01  g1978 ( .o(n7466), .a(n6571_1), .b(n5658) );
na02f01  g1979 ( .o(n7467), .a(n7466), .b(n5902) );
oa22f01  g1980 ( .o(n853), .a(n7467), .b(n5552_1), .c(n7465_1), .d(n7463) );
ao22f01  g1981 ( .o(n7469), .a(n5842), .b(net_9693), .c(n5841), .d(_net_131) );
na02f01  g1982 ( .o(n7470_1), .a(n5847), .b(net_9990) );
ao22f01  g1983 ( .o(n7471), .a(n5850), .b(net_9792), .c(n5849_1), .d(net_9891) );
na03f01  g1984 ( .o(n858), .a(n7471), .b(n7470_1), .c(n7469) );
na02f01  g1985 ( .o(n7473), .a(n7358), .b(net_256) );
na02f01  g1986 ( .o(n7474), .a(n7352), .b(net_9687) );
ao22f01  g1987 ( .o(n7475_1), .a(n7357), .b(_net_10120), .c(n7353), .d(x4359) );
na04f01  g1988 ( .o(n863), .a(n7475_1), .b(n7474), .c(n7473), .d(n7355_1) );
no02f01  g1989 ( .o(n7477), .a(n6886), .b(n5686) );
na02f01  g1990 ( .o(n7478), .a(n7477), .b(x6599) );
in01f01  g1991 ( .o(n7479), .a(n7477) );
na02f01  g1992 ( .o(n7480_1), .a(n7479), .b(x6599) );
oa22f01  g1993 ( .o(n868), .a(n7480_1), .b(n6778_1), .c(n7478), .d(n5561) );
in01f01  g1994 ( .o(n7482), .a(n6850) );
no03f01  g1995 ( .o(n7483), .a(n7482), .b(n6485), .c(n6504) );
no02f01  g1996 ( .o(n7484_1), .a(n6502), .b(n6504) );
na02f01  g1997 ( .o(n7485), .a(n7484_1), .b(n6853) );
no03f01  g1998 ( .o(n7486), .a(n7485), .b(n6505), .c(n6504) );
no03f01  g1999 ( .o(n7487), .a(n6861_1), .b(n6511), .c(n6504) );
na03f01  g2000 ( .o(n7488), .a(n6864), .b(_net_9243), .c(_net_9247) );
oa12f01  g2001 ( .o(n7489_1), .a(n7488), .b(n6477), .c(n6504) );
no04f01  g2002 ( .o(n7490), .a(n7489_1), .b(n7487), .c(n7486), .d(n7483) );
no02f01  g2003 ( .o(n7491), .a(n6467), .b(_net_9176) );
na02f01  g2004 ( .o(n7492), .a(n7491), .b(n6471) );
ao12f01  g2005 ( .o(n7493), .a(n6507_1), .b(n7492), .c(n7485) );
no03f01  g2006 ( .o(n7494_1), .a(n6474_1), .b(n6504), .c(n6463) );
ao22f01  g2007 ( .o(n7495), .a(n7484_1), .b(_net_9248), .c(n6494), .d(_net_9247) );
oa12f01  g2008 ( .o(n7496), .a(n7495), .b(n6499), .c(n6504) );
no03f01  g2009 ( .o(n7497), .a(n7496), .b(n7494_1), .c(n7493) );
ao12f01  g2010 ( .o(n873), .a(n6526_1), .b(n7497), .c(n7490) );
na02f01  g2011 ( .o(n7499_1), .a(net_115), .b(_net_9606) );
in01f01  g2012 ( .o(n7500), .a(_net_9606) );
in01f01  g2013 ( .o(n7501), .a(_net_9558) );
in01f01  g2014 ( .o(n7502), .a(_net_9636) );
no03f01  g2015 ( .o(n7503), .a(n5927), .b(n7502), .c(n7501) );
in01f01  g2016 ( .o(n7504_1), .a(n7503) );
ao12f01  g2017 ( .o(n7505), .a(_net_9558), .b(n5928), .c(_net_9636) );
in01f01  g2018 ( .o(n7506), .a(_net_9557) );
in01f01  g2019 ( .o(n7507), .a(_net_9635) );
no03f01  g2020 ( .o(n7508), .a(n5927), .b(n7507), .c(n7506) );
in01f01  g2021 ( .o(n7509_1), .a(n7508) );
oa12f01  g2022 ( .o(n7510), .a(n7504_1), .b(n7509_1), .c(n7505) );
ao12f01  g2023 ( .o(n7511), .a(_net_9557), .b(n5928), .c(_net_9635) );
no02f01  g2024 ( .o(n7512), .a(n7511), .b(n7505) );
na02f01  g2025 ( .o(n7513), .a(n5928), .b(net_9634) );
in01f01  g2026 ( .o(n7514_1), .a(n7513) );
in01f01  g2027 ( .o(n7515), .a(_net_9555) );
in01f01  g2028 ( .o(n7516), .a(_net_9300) );
oa22f01  g2029 ( .o(n7517), .a(n6026), .b(n7516), .c(n5923), .d(n5983_1) );
ao12f01  g2030 ( .o(n7518), .a(n7517), .b(n5928), .c(_net_9633) );
no02f01  g2031 ( .o(n7519_1), .a(n7518), .b(n7515) );
ao12f01  g2032 ( .o(n7520), .a(n7514_1), .b(n7519_1), .c(_net_9556) );
ao12f01  g2033 ( .o(n7521), .a(_net_9556), .b(n7519_1), .c(n7514_1) );
no02f01  g2034 ( .o(n7522), .a(n7514_1), .b(_net_9556) );
na02f01  g2035 ( .o(n7523), .a(n7518), .b(n7515) );
in01f01  g2036 ( .o(n7524_1), .a(n7523) );
no02f01  g2037 ( .o(n7525), .a(n7524_1), .b(n7522) );
in01f01  g2038 ( .o(n7526), .a(n7525) );
in01f01  g2039 ( .o(n7527), .a(net_9632) );
no02f01  g2040 ( .o(n7528), .a(n5927), .b(n7527) );
in01f01  g2041 ( .o(n7529_1), .a(_net_9299) );
no02f01  g2042 ( .o(n7530), .a(n6026), .b(n7529_1) );
no02f01  g2043 ( .o(n7531), .a(n5923), .b(n5990) );
no03f01  g2044 ( .o(n7532), .a(n7531), .b(n7530), .c(n7528) );
in01f01  g2045 ( .o(n7533), .a(n7532) );
in01f01  g2046 ( .o(n7534_1), .a(_net_9554) );
in01f01  g2047 ( .o(n7535), .a(_net_9553) );
in01f01  g2048 ( .o(n7536), .a(_net_9298) );
oa22f01  g2049 ( .o(n7537), .a(n6026), .b(n7536), .c(n5923), .d(n5989) );
ao12f01  g2050 ( .o(n7538_1), .a(n7537), .b(n5928), .c(net_9631) );
oa22f01  g2051 ( .o(n7539), .a(n7538_1), .b(n7535), .c(n7532), .d(n7534_1) );
oa12f01  g2052 ( .o(n7540), .a(n7539), .b(n7533), .c(_net_9554) );
oa22f01  g2053 ( .o(n7541), .a(n7540), .b(n7526), .c(n7521), .d(n7520) );
ao12f01  g2054 ( .o(n7542), .a(n7510), .b(n7541), .c(n7512) );
in01f01  g2055 ( .o(n7543_1), .a(n7542) );
na02f01  g2056 ( .o(n7544), .a(n5928), .b(_net_9629) );
in01f01  g2057 ( .o(n7545), .a(_net_9296) );
no02f01  g2058 ( .o(n7546), .a(n6026), .b(n7545) );
ao12f01  g2059 ( .o(n7547), .a(n7546), .b(n5924), .c(_net_173) );
na02f01  g2060 ( .o(n7548_1), .a(n7547), .b(n7544) );
na02f01  g2061 ( .o(n7549), .a(n7548_1), .b(_net_9551) );
in01f01  g2062 ( .o(n7550), .a(_net_9630) );
no02f01  g2063 ( .o(n7551), .a(n5927), .b(n7550) );
in01f01  g2064 ( .o(n7552_1), .a(_net_9297) );
no02f01  g2065 ( .o(n7553), .a(n6026), .b(n7552_1) );
in01f01  g2066 ( .o(n7554), .a(_net_174) );
no02f01  g2067 ( .o(n7555), .a(n5923), .b(n7554) );
no03f01  g2068 ( .o(n7556), .a(n7555), .b(n7553), .c(n7551) );
in01f01  g2069 ( .o(n7557_1), .a(n7556) );
na02f01  g2070 ( .o(n7558), .a(n7557_1), .b(_net_9552) );
no02f01  g2071 ( .o(n7559), .a(n7557_1), .b(_net_9552) );
ao22f01  g2072 ( .o(n7560), .a(n7559), .b(n7556), .c(n7558), .d(n7549) );
na02f01  g2073 ( .o(n7561), .a(n7560), .b(_net_9552) );
in01f01  g2074 ( .o(n7562_1), .a(n7559) );
in01f01  g2075 ( .o(n7563), .a(_net_9548) );
in01f01  g2076 ( .o(n7564), .a(net_9626) );
no02f01  g2077 ( .o(n7565), .a(n5927), .b(n7564) );
no02f01  g2078 ( .o(n7566_1), .a(n5923), .b(n7071) );
no03f01  g2079 ( .o(n7567), .a(n7566_1), .b(n7565), .c(n7074) );
in01f01  g2080 ( .o(n7568), .a(_net_9547) );
in01f01  g2081 ( .o(n7569), .a(net_9625) );
no02f01  g2082 ( .o(n7570), .a(n5927), .b(n7569) );
in01f01  g2083 ( .o(n7571_1), .a(_net_9292) );
no02f01  g2084 ( .o(n7572), .a(n6026), .b(n7571_1) );
in01f01  g2085 ( .o(n7573), .a(_net_169) );
no02f01  g2086 ( .o(n7574), .a(n5923), .b(n7573) );
no03f01  g2087 ( .o(n7575_1), .a(n7574), .b(n7572), .c(n7570) );
no02f01  g2088 ( .o(n7576), .a(n7575_1), .b(n7568) );
no02f01  g2089 ( .o(n7577), .a(n7567), .b(n7563) );
no02f01  g2090 ( .o(n7578), .a(n7577), .b(n7576) );
ao12f01  g2091 ( .o(n7579), .a(n7578), .b(n7567), .c(n7563) );
in01f01  g2092 ( .o(n7580_1), .a(n7579) );
in01f01  g2093 ( .o(n7581), .a(n7567) );
no02f01  g2094 ( .o(n7582), .a(n7581), .b(_net_9548) );
in01f01  g2095 ( .o(n7583), .a(n7582) );
na02f01  g2096 ( .o(n7584), .a(n7575_1), .b(n7568) );
in01f01  g2097 ( .o(n7585_1), .a(net_9624) );
no02f01  g2098 ( .o(n7586), .a(n5927), .b(n7585_1) );
oa22f01  g2099 ( .o(n7587), .a(n6026), .b(n6025), .c(n5923), .d(n5916) );
oa12f01  g2100 ( .o(n7588), .a(_net_9546), .b(n7587), .c(n7586) );
no03f01  g2101 ( .o(n7589), .a(n7587), .b(n7586), .c(_net_9546) );
in01f01  g2102 ( .o(n7590_1), .a(net_9623) );
no02f01  g2103 ( .o(n7591), .a(n5927), .b(n7590_1) );
in01f01  g2104 ( .o(n7592), .a(_net_167) );
in01f01  g2105 ( .o(n7593), .a(_net_9290) );
oa22f01  g2106 ( .o(n7594), .a(n6026), .b(n7593), .c(n5923), .d(n7592) );
oa12f01  g2107 ( .o(n7595_1), .a(net_9545), .b(n7594), .c(n7591) );
oa12f01  g2108 ( .o(n7596), .a(n7588), .b(n7595_1), .c(n7589) );
na03f01  g2109 ( .o(n7597), .a(n7596), .b(n7584), .c(n7583) );
no02f01  g2110 ( .o(n7598), .a(n7548_1), .b(_net_9551) );
na02f01  g2111 ( .o(n7599), .a(n5928), .b(_net_9628) );
na02f01  g2112 ( .o(n7600_1), .a(n5924), .b(_net_172) );
na03f01  g2113 ( .o(n7601), .a(n5925), .b(n5923), .c(_net_9295) );
na03f01  g2114 ( .o(n7602), .a(n7601), .b(n7600_1), .c(n7599) );
no02f01  g2115 ( .o(n7603), .a(n7602), .b(_net_9550) );
na02f01  g2116 ( .o(n7604), .a(n5928), .b(_net_9627) );
in01f01  g2117 ( .o(n7605_1), .a(_net_9294) );
no02f01  g2118 ( .o(n7606), .a(n6026), .b(n7605_1) );
ao12f01  g2119 ( .o(n7607), .a(n7606), .b(n5924), .c(_net_171) );
na02f01  g2120 ( .o(n7608), .a(n7607), .b(n7604) );
no02f01  g2121 ( .o(n7609_1), .a(n7608), .b(net_9549) );
no03f01  g2122 ( .o(n7610), .a(n7609_1), .b(n7603), .c(n7598) );
in01f01  g2123 ( .o(n7611), .a(n7610) );
ao12f01  g2124 ( .o(n7612), .a(n7611), .b(n7597), .c(n7580_1) );
na02f01  g2125 ( .o(n7613_1), .a(n7602), .b(_net_9550) );
na02f01  g2126 ( .o(n7614), .a(n7613_1), .b(n7603) );
na02f01  g2127 ( .o(n7615), .a(n7608), .b(net_9549) );
ao12f01  g2128 ( .o(n7616), .a(n7598), .b(n7615), .c(n7613_1) );
ao12f01  g2129 ( .o(n7617_1), .a(n7560), .b(n7616), .c(n7614) );
in01f01  g2130 ( .o(n7618), .a(n7617_1) );
oa12f01  g2131 ( .o(n7619), .a(n7562_1), .b(n7618), .c(n7612) );
na02f01  g2132 ( .o(n7620), .a(n7538_1), .b(n7535) );
oa12f01  g2133 ( .o(n7621_1), .a(n7620), .b(n7533), .c(_net_9554) );
no02f01  g2134 ( .o(n7622), .a(n7621_1), .b(n7526) );
in01f01  g2135 ( .o(n7623), .a(n7622) );
ao12f01  g2136 ( .o(n7624), .a(n7623), .b(n7619), .c(n7561) );
in01f01  g2137 ( .o(n7625), .a(net_9559) );
in01f01  g2138 ( .o(n7626_1), .a(n7512) );
no02f01  g2139 ( .o(n7627), .a(n7626_1), .b(n7625) );
ao22f01  g2140 ( .o(n7628), .a(n7627), .b(n7624), .c(n7543_1), .d(net_9559) );
no02f01  g2141 ( .o(n7629), .a(n7628), .b(net_9560) );
in01f01  g2142 ( .o(n7630), .a(net_9560) );
in01f01  g2143 ( .o(n7631_1), .a(n7561) );
na02f01  g2144 ( .o(n7632), .a(n7596), .b(n7584) );
no02f01  g2145 ( .o(n7633), .a(n7632), .b(n7582) );
oa12f01  g2146 ( .o(n7634), .a(n7610), .b(n7633), .c(n7579) );
ao12f01  g2147 ( .o(n7635), .a(n7559), .b(n7617_1), .c(n7634) );
oa12f01  g2148 ( .o(n7636_1), .a(n7622), .b(n7635), .c(n7631_1) );
in01f01  g2149 ( .o(n7637), .a(n7627) );
oa22f01  g2150 ( .o(n7638), .a(n7637), .b(n7636_1), .c(n7542), .d(n7625) );
no02f01  g2151 ( .o(n7639), .a(n7638), .b(n7630) );
oa12f01  g2152 ( .o(n7640_1), .a(n7500), .b(n7639), .c(n7629) );
na02f01  g2153 ( .o(n878), .a(n7640_1), .b(n7499_1) );
ao22f01  g2154 ( .o(n7642), .a(n6602), .b(net_10005), .c(n6555), .d(net_9973) );
ao22f01  g2155 ( .o(n7643), .a(n6582), .b(net_9906), .c(n6573), .d(net_9874) );
ao22f01  g2156 ( .o(n7644), .a(n6585), .b(net_9708), .c(n6577), .d(net_9676) );
ao22f01  g2157 ( .o(n7645_1), .a(n6584_1), .b(net_9775), .c(n6580), .d(net_9807) );
na04f01  g2158 ( .o(n883), .a(n7645_1), .b(n7644), .c(n7643), .d(n7642) );
na02f01  g2159 ( .o(n7647), .a(n6693), .b(n6692) );
na02f01  g2160 ( .o(n7648), .a(n7647), .b(n6695) );
oa22f01  g2161 ( .o(n888), .a(n7648), .b(n6688), .c(n6685), .d(n6692) );
in01f01  g2162 ( .o(n7650_1), .a(net_9208) );
in01f01  g2163 ( .o(n7651), .a(_net_9207) );
no02f01  g2164 ( .o(n7652), .a(n6704_1), .b(n7651) );
in01f01  g2165 ( .o(n7653), .a(n7652) );
no02f01  g2166 ( .o(n7654), .a(n7653), .b(n7650_1) );
oa12f01  g2167 ( .o(n7655_1), .a(n6687), .b(n7652), .c(net_9208) );
oa22f01  g2168 ( .o(n893), .a(n7655_1), .b(n7654), .c(n6685), .d(n7650_1) );
ao12f01  g2169 ( .o(n7657), .a(n5658), .b(n6532), .c(net_245) );
ao22f01  g2170 ( .o(n7658), .a(n6535), .b(x5225), .c(n6534), .d(net_10005) );
na02f01  g2171 ( .o(n898), .a(n7658), .b(n7657) );
in01f01  g2172 ( .o(n7660_1), .a(n6544) );
no02f01  g2173 ( .o(n7661), .a(n6543), .b(net_9616) );
no03f01  g2174 ( .o(n903), .a(n7661), .b(n7660_1), .c(net_9613) );
no02f01  g2175 ( .o(n7663), .a(_net_10433), .b(_net_10434) );
in01f01  g2176 ( .o(n7664), .a(n7663) );
ao12f01  g2177 ( .o(n7665_1), .a(_net_10431), .b(_net_10430), .c(_net_10429) );
in01f01  g2178 ( .o(n7666), .a(n7665_1) );
no02f01  g2179 ( .o(n7667), .a(n7666), .b(_net_10432) );
in01f01  g2180 ( .o(n7668), .a(n7667) );
no02f01  g2181 ( .o(n7669), .a(n7668), .b(n7664) );
in01f01  g2182 ( .o(n7670_1), .a(n7669) );
no02f01  g2183 ( .o(n7671), .a(n7670_1), .b(_net_10435) );
in01f01  g2184 ( .o(n7672), .a(n7671) );
no02f01  g2185 ( .o(n7673), .a(n7672), .b(_net_10436) );
in01f01  g2186 ( .o(n7674), .a(n7673) );
no02f01  g2187 ( .o(n7675_1), .a(n7674), .b(_net_10437) );
in01f01  g2188 ( .o(n7676), .a(n7675_1) );
no02f01  g2189 ( .o(n7677), .a(n7676), .b(_net_10438) );
in01f01  g2190 ( .o(n7678), .a(n7677) );
na02f01  g2191 ( .o(n7679), .a(n7676), .b(_net_10438) );
na02f01  g2192 ( .o(n908), .a(n7679), .b(n7678) );
no02f01  g2193 ( .o(n7681), .a(n6904), .b(_net_10248) );
no02f01  g2194 ( .o(n7682), .a(n6783), .b(n7681) );
oa12f01  g2195 ( .o(n7683), .a(n7682), .b(n6793), .c(n6782_1) );
no03f01  g2196 ( .o(n7684), .a(n7682), .b(n6793), .c(n6782_1) );
no02f01  g2197 ( .o(n7685_1), .a(n7684), .b(n6933) );
na02f01  g2198 ( .o(n7686), .a(n7685_1), .b(n7683) );
no02f01  g2199 ( .o(n7687), .a(n6832), .b(_net_10248) );
no02f01  g2200 ( .o(n7688), .a(n7687), .b(n6834) );
ao22f01  g2201 ( .o(n7689), .a(n7688), .b(n6175), .c(n6168), .d(_net_10248) );
na02f01  g2202 ( .o(n913), .a(n7689), .b(n7686) );
in01f01  g2203 ( .o(n7691), .a(_net_10203) );
ao12f01  g2204 ( .o(n7692), .a(n5658), .b(n6887), .c(x5901) );
oa12f01  g2205 ( .o(n922), .a(n7692), .b(n6885_1), .c(n7691) );
ao22f01  g2206 ( .o(n7694), .a(n5842), .b(net_9684), .c(n5841), .d(_net_122) );
na02f01  g2207 ( .o(n7695_1), .a(n5847), .b(net_9981) );
ao22f01  g2208 ( .o(n7696), .a(n5850), .b(net_9783), .c(n5849_1), .d(net_9882) );
na03f01  g2209 ( .o(n927), .a(n7696), .b(n7695_1), .c(n7694) );
in01f01  g2210 ( .o(n7698), .a(_net_9232) );
na03f01  g2211 ( .o(n7699), .a(n6486), .b(n6484_1), .c(_net_9237) );
na03f01  g2212 ( .o(n7700_1), .a(n6516), .b(n6513), .c(_net_9236) );
na03f01  g2213 ( .o(n7701), .a(n7700_1), .b(n7699), .c(n6520) );
no02f01  g2214 ( .o(n7702), .a(n7701), .b(n6515) );
na02f01  g2215 ( .o(n7703), .a(n7702), .b(n7698) );
na02f01  g2216 ( .o(n7704_1), .a(net_9228), .b(net_9229) );
in01f01  g2217 ( .o(n7705), .a(n7704_1) );
no02f01  g2218 ( .o(n7706), .a(net_9228), .b(net_9229) );
no03f01  g2219 ( .o(n936), .a(n7706), .b(n7705), .c(n7703) );
in01f01  g2220 ( .o(n7708), .a(net_9257) );
na02f01  g2221 ( .o(n7709_1), .a(n6349), .b(n6290) );
oa22f01  g2222 ( .o(n949), .a(n7709_1), .b(n6348), .c(n6349), .d(n7708) );
oa22f01  g2223 ( .o(n954), .a(n7480_1), .b(n6776), .c(n7478), .d(n5649) );
na02f01  g2224 ( .o(n7712), .a(n6038), .b(net_251) );
na02f01  g2225 ( .o(n7713), .a(n6037_1), .b(net_9880) );
ao22f01  g2226 ( .o(n7714_1), .a(n6044), .b(x4781), .c(n6042_1), .d(_net_10325) );
na04f01  g2227 ( .o(n963), .a(n7714_1), .b(n7713), .c(n7712), .d(n6040) );
no02f01  g2228 ( .o(n7716), .a(n6545), .b(net_9618) );
no03f01  g2229 ( .o(n973), .a(n7716), .b(n6547), .c(net_9613) );
in01f01  g2230 ( .o(n7718), .a(x3632) );
no02f01  g2231 ( .o(n982), .a(n7718), .b(n5658) );
in01f01  g2232 ( .o(n7720), .a(_net_9562) );
na02f01  g2233 ( .o(n7721), .a(n6009_1), .b(_net_9564) );
na03f01  g2234 ( .o(n7722), .a(n5935_1), .b(n5929), .c(net_9570) );
in01f01  g2235 ( .o(n7723), .a(_net_187) );
no02f01  g2236 ( .o(n7724_1), .a(_net_188), .b(n7723) );
in01f01  g2237 ( .o(n7725), .a(n7724_1) );
no02f01  g2238 ( .o(n7726), .a(n7725), .b(_net_8833) );
no03f01  g2239 ( .o(n7727), .a(_net_8834), .b(n5918), .c(_net_187) );
oa12f01  g2240 ( .o(n7728), .a(n5922), .b(n7727), .c(n7726) );
na04f01  g2241 ( .o(n997), .a(n7728), .b(n7722), .c(n7721), .d(n7720) );
in01f01  g2242 ( .o(n7730), .a(_net_9346) );
in01f01  g2243 ( .o(n7731), .a(net_9155) );
in01f01  g2244 ( .o(n7732), .a(net_9151) );
in01f01  g2245 ( .o(n7733), .a(_net_9161) );
no02f01  g2246 ( .o(n7734_1), .a(n7733), .b(n7732) );
no03f01  g2247 ( .o(n7735), .a(_net_9355), .b(_net_9356), .c(_net_9354) );
na03f01  g2248 ( .o(n7736), .a(n7735), .b(n7734_1), .c(x6599) );
ao12f01  g2249 ( .o(n7737), .a(n5658), .b(n7735), .c(n7734_1) );
in01f01  g2250 ( .o(n7738_1), .a(n7737) );
oa22f01  g2251 ( .o(n1002), .a(n7738_1), .b(n7730), .c(n7736), .d(n7731) );
in01f01  g2252 ( .o(n7740), .a(net_9175) );
in01f01  g2253 ( .o(n7741), .a(_net_9173) );
in01f01  g2254 ( .o(n7742), .a(net_9174) );
no02f01  g2255 ( .o(n7743_1), .a(n7742), .b(n7741) );
in01f01  g2256 ( .o(n7744), .a(n7743_1) );
no02f01  g2257 ( .o(n7745), .a(n7744), .b(net_9175) );
no02f01  g2258 ( .o(n7746), .a(n7743_1), .b(n7740) );
no02f01  g2259 ( .o(n7747), .a(n6483), .b(_net_9176) );
ao22f01  g2260 ( .o(n7748_1), .a(n7747), .b(_net_9247), .c(n7491), .d(_net_9246) );
no02f01  g2261 ( .o(n5656), .a(n7748_1), .b(_net_9245) );
oa12f01  g2262 ( .o(n7750), .a(n5656), .b(n7746), .c(n7745) );
na02f01  g2263 ( .o(n7751), .a(n7748_1), .b(n6475) );
oa12f01  g2264 ( .o(n1007), .a(n7750), .b(n7751), .c(n7740) );
in01f01  g2265 ( .o(n7753_1), .a(net_217) );
in01f01  g2266 ( .o(n7754), .a(_net_9272) );
na02f01  g2267 ( .o(n7755), .a(n7754), .b(x6599) );
na02f01  g2268 ( .o(n7756), .a(_net_9272), .b(x6599) );
oa22f01  g2269 ( .o(n1012), .a(n7756), .b(n5779), .c(n7755), .d(n7753_1) );
ao12f01  g2270 ( .o(n7758_1), .a(n5658), .b(n6532), .c(_net_234) );
ao22f01  g2271 ( .o(n7759), .a(n6535), .b(x5901), .c(n6534), .d(net_9994) );
na02f01  g2272 ( .o(n1017), .a(n7759), .b(n7758_1) );
in01f01  g2273 ( .o(n7761), .a(_net_10122) );
no02f01  g2274 ( .o(n7762), .a(n7761), .b(_net_10160) );
in01f01  g2275 ( .o(n7763_1), .a(_net_10160) );
no02f01  g2276 ( .o(n7764), .a(_net_10122), .b(n7763_1) );
in01f01  g2277 ( .o(n7765), .a(_net_10159) );
no02f01  g2278 ( .o(n7766), .a(_net_10121), .b(n7765) );
in01f01  g2279 ( .o(n7767), .a(_net_10156) );
no02f01  g2280 ( .o(n7768_1), .a(_net_10118), .b(n7767) );
in01f01  g2281 ( .o(n7769), .a(_net_10155) );
no02f01  g2282 ( .o(n7770), .a(n7769), .b(_net_10117) );
in01f01  g2283 ( .o(n7771), .a(_net_10117) );
in01f01  g2284 ( .o(n7772), .a(_net_10116) );
no02f01  g2285 ( .o(n7773_1), .a(_net_10154), .b(n7772) );
in01f01  g2286 ( .o(n7774), .a(n7773_1) );
oa12f01  g2287 ( .o(n7775), .a(n7771), .b(n7774), .c(_net_10155) );
oa12f01  g2288 ( .o(n7776), .a(_net_10155), .b(n7774), .c(n7771) );
na02f01  g2289 ( .o(n7777), .a(n7776), .b(n7775) );
in01f01  g2290 ( .o(n7778_1), .a(_net_10154) );
no02f01  g2291 ( .o(n7779), .a(n7778_1), .b(_net_10116) );
in01f01  g2292 ( .o(n7780), .a(_net_10115) );
no02f01  g2293 ( .o(n7781), .a(_net_10153), .b(n7780) );
in01f01  g2294 ( .o(n7782_1), .a(_net_10152) );
no02f01  g2295 ( .o(n7783), .a(n7782_1), .b(_net_10114) );
in01f01  g2296 ( .o(n7784), .a(n7783) );
in01f01  g2297 ( .o(n7785), .a(_net_10153) );
no02f01  g2298 ( .o(n7786), .a(n7785), .b(_net_10115) );
in01f01  g2299 ( .o(n7787_1), .a(n7786) );
ao12f01  g2300 ( .o(n7788), .a(n7781), .b(n7787_1), .c(n7784) );
no02f01  g2301 ( .o(n7789), .a(n7788), .b(n7779) );
in01f01  g2302 ( .o(n7790), .a(n7789) );
oa12f01  g2303 ( .o(n7791), .a(n7777), .b(n7790), .c(n7770) );
in01f01  g2304 ( .o(n7792_1), .a(n7791) );
no02f01  g2305 ( .o(n7793), .a(n7792_1), .b(n7768_1) );
in01f01  g2306 ( .o(n7794), .a(_net_10158) );
no02f01  g2307 ( .o(n7795), .a(_net_10120), .b(n7794) );
in01f01  g2308 ( .o(n7796_1), .a(n7795) );
in01f01  g2309 ( .o(n7797), .a(_net_10157) );
no02f01  g2310 ( .o(n7798), .a(n7797), .b(_net_10119) );
in01f01  g2311 ( .o(n7799), .a(n7798) );
na03f01  g2312 ( .o(n7800), .a(n7799), .b(n7796_1), .c(n7793) );
in01f01  g2313 ( .o(n7801_1), .a(_net_10119) );
no02f01  g2314 ( .o(n7802), .a(_net_10157), .b(n7801_1) );
in01f01  g2315 ( .o(n7803), .a(_net_10118) );
no02f01  g2316 ( .o(n7804), .a(n7803), .b(_net_10156) );
ao12f01  g2317 ( .o(n7805), .a(n7802), .b(n7804), .c(n7799) );
no02f01  g2318 ( .o(n7806_1), .a(n7805), .b(n7795) );
in01f01  g2319 ( .o(n7807), .a(_net_10121) );
in01f01  g2320 ( .o(n7808), .a(_net_10120) );
no02f01  g2321 ( .o(n7809), .a(n7808), .b(_net_10158) );
no02f01  g2322 ( .o(n7810), .a(n7807), .b(_net_10159) );
no02f01  g2323 ( .o(n7811_1), .a(n7810), .b(n7809) );
ao12f01  g2324 ( .o(n7812), .a(n7811_1), .b(n7766), .c(n7807) );
no02f01  g2325 ( .o(n7813), .a(n7812), .b(n7806_1) );
ao12f01  g2326 ( .o(n7814), .a(n7766), .b(n7813), .c(n7800) );
na02f01  g2327 ( .o(n7815), .a(n7812), .b(n7765) );
in01f01  g2328 ( .o(n7816_1), .a(n7815) );
no02f01  g2329 ( .o(n7817), .a(n7816_1), .b(n7814) );
no02f01  g2330 ( .o(n7818), .a(n7817), .b(n7764) );
no02f01  g2331 ( .o(n7819), .a(n7818), .b(n7762) );
in01f01  g2332 ( .o(n7820), .a(_net_10161) );
no02f01  g2333 ( .o(n7821_1), .a(n7820), .b(_net_10123) );
in01f01  g2334 ( .o(n7822), .a(_net_10123) );
no02f01  g2335 ( .o(n7823), .a(_net_10161), .b(n7822) );
no02f01  g2336 ( .o(n7824), .a(n7823), .b(n7821_1) );
na02f01  g2337 ( .o(n7825), .a(n7824), .b(n7819) );
in01f01  g2338 ( .o(n7826_1), .a(n7824) );
oa12f01  g2339 ( .o(n7827), .a(n7826_1), .b(n7818), .c(n7762) );
na02f01  g2340 ( .o(n1022), .a(n7827), .b(n7825) );
no03f01  g2341 ( .o(n7829), .a(n6643), .b(n6642), .c(n6638) );
no02f01  g2342 ( .o(n7830_1), .a(n6644_1), .b(n6615) );
na02f01  g2343 ( .o(n7831), .a(n7830_1), .b(n7829) );
in01f01  g2344 ( .o(n7832), .a(n7829) );
in01f01  g2345 ( .o(n7833), .a(n7830_1) );
na02f01  g2346 ( .o(n7834_1), .a(n7833), .b(n7832) );
na02f01  g2347 ( .o(n1027), .a(n7834_1), .b(n7831) );
ao22f01  g2348 ( .o(n7836), .a(n5842), .b(net_9681), .c(n5841), .d(_net_119) );
na02f01  g2349 ( .o(n7837), .a(n5847), .b(net_9978) );
ao22f01  g2350 ( .o(n7838), .a(n5850), .b(net_9780), .c(n5849_1), .d(net_9879) );
na03f01  g2351 ( .o(n1037), .a(n7838), .b(n7837), .c(n7836) );
no02f01  g2352 ( .o(n7840), .a(n6886), .b(n5660) );
in01f01  g2353 ( .o(n7841), .a(net_10280) );
no02f01  g2354 ( .o(n7842), .a(n5675), .b(n7841) );
in01f01  g2355 ( .o(n7843_1), .a(n7842) );
no03f01  g2356 ( .o(n7844), .a(n7843_1), .b(n7840), .c(n5658) );
ao12f01  g2357 ( .o(n7845), .a(n5658), .b(n7844), .c(net_256) );
no03f01  g2358 ( .o(n7846), .a(n7842), .b(n7840), .c(n5658) );
no03f01  g2359 ( .o(n7847), .a(n6886), .b(n5660), .c(n5658) );
ao22f01  g2360 ( .o(n7848_1), .a(n7847), .b(x4359), .c(n7846), .d(net_9818) );
na02f01  g2361 ( .o(n1042), .a(n7848_1), .b(n7845) );
no02f01  g2362 ( .o(n7850), .a(n6513), .b(n6479_1) );
oa12f01  g2363 ( .o(n7851), .a(n6516), .b(n7850), .c(n6674_1) );
in01f01  g2364 ( .o(n7852), .a(_net_9248) );
na02f01  g2365 ( .o(n7853_1), .a(n6471), .b(_net_9237) );
no02f01  g2366 ( .o(n7854), .a(n7853_1), .b(n7852) );
na03f01  g2367 ( .o(n7855), .a(n6864), .b(_net_9243), .c(_net_9237) );
oa12f01  g2368 ( .o(n7856), .a(n7855), .b(n6477), .c(n6479_1) );
no02f01  g2369 ( .o(n7857_1), .a(n7856), .b(n7854) );
oa12f01  g2370 ( .o(n7858), .a(n7857_1), .b(n7851), .c(n6511) );
ao12f01  g2371 ( .o(n7859), .a(n7858), .b(n6850), .c(n6486) );
no03f01  g2372 ( .o(n7860), .a(n6474_1), .b(n6479_1), .c(n6463) );
ao12f01  g2373 ( .o(n7861), .a(n6479_1), .b(n6499), .c(n6493_1) );
in01f01  g2374 ( .o(n7862_1), .a(n6506) );
in01f01  g2375 ( .o(n7863), .a(n6508) );
ao12f01  g2376 ( .o(n7864), .a(n7853_1), .b(n7863), .c(n7862_1) );
no03f01  g2377 ( .o(n7865), .a(n7864), .b(n7861), .c(n7860) );
ao12f01  g2378 ( .o(n1047), .a(n6526_1), .b(n7865), .c(n7859) );
ao12f01  g2379 ( .o(n7867), .a(n5658), .b(n5678), .c(net_249) );
ao22f01  g2380 ( .o(n7868), .a(n5681_1), .b(x4937), .c(n5680), .d(net_9712) );
na02f01  g2381 ( .o(n1052), .a(n7868), .b(n7867) );
no02f01  g2382 ( .o(n7870), .a(n7404), .b(n7390) );
in01f01  g2383 ( .o(n7871_1), .a(_net_10028) );
no02f01  g2384 ( .o(n7872), .a(n7871_1), .b(n7433) );
no02f01  g2385 ( .o(n7873), .a(n7872), .b(n7386) );
in01f01  g2386 ( .o(n7874), .a(n7873) );
in01f01  g2387 ( .o(n7875), .a(n7431) );
ao12f01  g2388 ( .o(n7876_1), .a(n7875), .b(n7874), .c(n7870) );
oa12f01  g2389 ( .o(n7877), .a(n7876_1), .b(n7874), .c(n7870) );
oa12f01  g2390 ( .o(n7878), .a(_net_10470), .b(n7435), .c(_net_10469) );
ao12f01  g2391 ( .o(n7879), .a(n7451_1), .b(n7878), .c(n7437) );
ao12f01  g2392 ( .o(n7880), .a(n7879), .b(n7453), .c(_net_10470) );
na02f01  g2393 ( .o(n1057), .a(n7880), .b(n7877) );
in01f01  g2394 ( .o(n7882), .a(_net_9325) );
no02f01  g2395 ( .o(n7883), .a(n7732), .b(_net_9351) );
in01f01  g2396 ( .o(n7884), .a(_net_9356) );
in01f01  g2397 ( .o(n7885_1), .a(n7734_1) );
no02f01  g2398 ( .o(n7886), .a(n7885_1), .b(_net_9160) );
in01f01  g2399 ( .o(n7887), .a(n7886) );
in01f01  g2400 ( .o(n7888), .a(_net_9160) );
in01f01  g2401 ( .o(n7889_1), .a(_net_9354) );
in01f01  g2402 ( .o(n7890), .a(_net_9344) );
no02f01  g2403 ( .o(n7891), .a(_net_9343), .b(n7890) );
in01f01  g2404 ( .o(n7892), .a(n7891) );
no02f01  g2405 ( .o(n7893_1), .a(_net_9345), .b(_net_9346) );
in01f01  g2406 ( .o(n7894), .a(n7893_1) );
no02f01  g2407 ( .o(n7895), .a(n7894), .b(n7892) );
ao12f01  g2408 ( .o(n7896), .a(n7889_1), .b(n7895), .c(n7888) );
no02f01  g2409 ( .o(n7897), .a(n6454), .b(n7890) );
in01f01  g2410 ( .o(n7898_1), .a(n7897) );
no02f01  g2411 ( .o(n7899), .a(n7898_1), .b(n7894) );
no02f01  g2412 ( .o(n7900), .a(n6457), .b(n7730) );
in01f01  g2413 ( .o(n7901), .a(n7900) );
no02f01  g2414 ( .o(n7902_1), .a(n7901), .b(n7898_1) );
no02f01  g2415 ( .o(n7903), .a(_net_9345), .b(n7730) );
in01f01  g2416 ( .o(n7904), .a(n7903) );
no02f01  g2417 ( .o(n7905), .a(n7904), .b(n7898_1) );
no02f01  g2418 ( .o(n7906_1), .a(n7898_1), .b(n6459) );
no04f01  g2419 ( .o(n7907), .a(n7906_1), .b(n7905), .c(n7902_1), .d(n7899) );
no02f01  g2420 ( .o(n7908), .a(n7907), .b(n7887) );
no02f01  g2421 ( .o(n2439), .a(n7901), .b(n6456_1) );
in01f01  g2422 ( .o(n7910), .a(n2439) );
no02f01  g2423 ( .o(n2740), .a(n7904), .b(n6456_1) );
no02f01  g2424 ( .o(n3455), .a(n7894), .b(n6456_1) );
no02f01  g2425 ( .o(n7913), .a(n3455), .b(n2740) );
na02f01  g2426 ( .o(n7914), .a(n7913), .b(n7910) );
in01f01  g2427 ( .o(n7915), .a(n7914) );
no02f01  g2428 ( .o(n7916_1), .a(_net_9343), .b(_net_9344) );
in01f01  g2429 ( .o(n7917), .a(n7916_1) );
no02f01  g2430 ( .o(n8021), .a(n7917), .b(n6459) );
no02f01  g2431 ( .o(n7919), .a(n8021), .b(n6460_1) );
na02f01  g2432 ( .o(n7920), .a(n7919), .b(n7915) );
na02f01  g2433 ( .o(n7921_1), .a(n7920), .b(n7886) );
na03f01  g2434 ( .o(n7922), .a(n7921_1), .b(n7908), .c(n7896) );
oa12f01  g2435 ( .o(n7923), .a(n7922), .b(n7887), .c(n7884) );
no02f01  g2436 ( .o(n7924), .a(n7923), .b(n7883) );
in01f01  g2437 ( .o(n7925_1), .a(n7924) );
ao12f01  g2438 ( .o(n7926), .a(n7883), .b(n7923), .c(_net_9317) );
oa12f01  g2439 ( .o(n1062), .a(n7926), .b(n7925_1), .c(n7882) );
ao12f01  g2440 ( .o(n7928), .a(n5658), .b(n5678), .c(_net_231) );
ao22f01  g2441 ( .o(n7929), .a(n5681_1), .b(x6102), .c(n5680), .d(net_9694) );
na02f01  g2442 ( .o(n1067), .a(n7929), .b(n7928) );
in01f01  g2443 ( .o(n7931), .a(n6885_1) );
na04f01  g2444 ( .o(n7932), .a(n7931), .b(_net_133), .c(net_10280), .d(n6031) );
na03f01  g2445 ( .o(n7933), .a(n7931), .b(net_10280), .c(_net_132) );
no02f01  g2446 ( .o(n7934), .a(n6887), .b(n5658) );
na03f01  g2447 ( .o(n7935_1), .a(n7934), .b(n7933), .c(n7932) );
in01f01  g2448 ( .o(n7936), .a(n7935_1) );
no02f01  g2449 ( .o(n7937), .a(n7936), .b(n7932) );
na02f01  g2450 ( .o(n7938), .a(n7937), .b(net_244) );
na02f01  g2451 ( .o(n7939), .a(n7935_1), .b(n5658) );
na02f01  g2452 ( .o(n7940_1), .a(n7936), .b(net_9774) );
in01f01  g2453 ( .o(n7941), .a(n6887) );
no02f01  g2454 ( .o(n7942), .a(n7936), .b(n7941) );
no02f01  g2455 ( .o(n7943), .a(n7936), .b(n7933) );
ao22f01  g2456 ( .o(n7944), .a(n7943), .b(_net_10213), .c(n7942), .d(x5289) );
na04f01  g2457 ( .o(n1072), .a(n7944), .b(n7940_1), .c(n7939), .d(n7938) );
na02f01  g2458 ( .o(n7946), .a(n7358), .b(net_247) );
na02f01  g2459 ( .o(n7947), .a(n7352), .b(net_9678) );
ao22f01  g2460 ( .o(n7948), .a(n7357), .b(_net_10111), .c(n7353), .d(x5077) );
na04f01  g2461 ( .o(n1077), .a(n7948), .b(n7947), .c(n7946), .d(n7355_1) );
ao22f01  g2462 ( .o(n7950_1), .a(n5842), .b(net_9701), .c(n5841), .d(net_141) );
na02f01  g2463 ( .o(n7951), .a(n5847), .b(net_9998) );
ao22f01  g2464 ( .o(n7952), .a(n5850), .b(net_9800), .c(n5849_1), .d(net_9899) );
na03f01  g2465 ( .o(n1082), .a(n7952), .b(n7951), .c(n7950_1) );
in01f01  g2466 ( .o(n7954_1), .a(net_10179) );
no02f01  g2467 ( .o(n7955), .a(n7464), .b(n6158) );
na02f01  g2468 ( .o(n7956), .a(n7466), .b(n5671_1) );
oa22f01  g2469 ( .o(n1087), .a(n7956), .b(n5637), .c(n7955), .d(n7954_1) );
in01f01  g2470 ( .o(n7958), .a(n2740) );
no02f01  g2471 ( .o(n7959), .a(n7958), .b(n5931_1) );
oa12f01  g2472 ( .o(n7960), .a(_net_9565), .b(n7959), .c(_net_9562) );
na03f01  g2473 ( .o(n7961), .a(n3455), .b(n5921_1), .c(_net_9562) );
na02f01  g2474 ( .o(n7962_1), .a(n7961), .b(n7728) );
in01f01  g2475 ( .o(n7963), .a(n7962_1) );
na02f01  g2476 ( .o(n7964), .a(n7963), .b(n7960) );
in01f01  g2477 ( .o(n7965), .a(_net_184) );
no02f01  g2478 ( .o(n7966), .a(_net_183), .b(n7965) );
in01f01  g2479 ( .o(n7967_1), .a(n7966) );
na02f01  g2480 ( .o(n7968), .a(n8021), .b(net_313) );
na02f01  g2481 ( .o(n7969), .a(n7968), .b(n7967_1) );
in01f01  g2482 ( .o(n7970), .a(_net_9573) );
ao12f01  g2483 ( .o(n7971), .a(n7970), .b(_net_183), .c(n7965) );
na02f01  g2484 ( .o(n7972_1), .a(n7971), .b(n6461) );
no03f01  g2485 ( .o(n7973), .a(n7972_1), .b(n7969), .c(n7964) );
no02f01  g2486 ( .o(n7974), .a(n7959), .b(n7724_1) );
in01f01  g2487 ( .o(n7975), .a(n7974) );
na03f01  g2488 ( .o(n7976), .a(n7975), .b(n7973), .c(_net_9637) );
na02f01  g2489 ( .o(n7977_1), .a(n7976), .b(n5855) );
in01f01  g2490 ( .o(n7978), .a(n7977_1) );
in01f01  g2491 ( .o(n7979), .a(_net_9536) );
no02f01  g2492 ( .o(n7980), .a(n5489), .b(n7979) );
no04f01  g2493 ( .o(n7981), .a(_net_9521), .b(net_9526), .c(_net_9520), .d(_net_9519) );
no04f01  g2494 ( .o(n7982_1), .a(net_9529), .b(net_9527), .c(net_9528), .d(_net_9518) );
na02f01  g2495 ( .o(n7983), .a(n7982_1), .b(n7981) );
no04f01  g2496 ( .o(n7984), .a(net_9523), .b(net_9522), .c(net_9524), .d(net_9525) );
in01f01  g2497 ( .o(n7985), .a(n7984) );
no02f01  g2498 ( .o(n7986), .a(_net_9517), .b(_net_9516) );
in01f01  g2499 ( .o(n7987_1), .a(n7986) );
no03f01  g2500 ( .o(n3300), .a(n7987_1), .b(n7985), .c(n7983) );
in01f01  g2501 ( .o(n7989), .a(n3300) );
ao12f01  g2502 ( .o(n7990), .a(n7980), .b(n7989), .c(n6132) );
no02f01  g2503 ( .o(n7991), .a(n7978), .b(n5658) );
na02f01  g2504 ( .o(n7992_1), .a(n6020), .b(n6625) );
oa12f01  g2505 ( .o(n3364), .a(n7992_1), .b(n6020), .c(n7573) );
na02f01  g2506 ( .o(n7994), .a(n3364), .b(n7991) );
no02f01  g2507 ( .o(n7995), .a(n7987_1), .b(_net_9518) );
in01f01  g2508 ( .o(n7996_1), .a(n7995) );
na02f01  g2509 ( .o(n7997), .a(n7987_1), .b(_net_9518) );
no03f01  g2510 ( .o(n7998), .a(n7990), .b(n7977_1), .c(n5658) );
in01f01  g2511 ( .o(n7999), .a(n7998) );
ao12f01  g2512 ( .o(n8000), .a(n7999), .b(n7997), .c(n7996_1) );
in01f01  g2513 ( .o(n8001_1), .a(_net_9518) );
na03f01  g2514 ( .o(n8002), .a(n7990), .b(n7978), .c(x6599) );
oa12f01  g2515 ( .o(n8003), .a(x6599), .b(n8002), .c(n8001_1) );
no02f01  g2516 ( .o(n8004), .a(n8003), .b(n8000) );
na02f01  g2517 ( .o(n1092), .a(n8004), .b(n7994) );
ao22f01  g2518 ( .o(n8006_1), .a(n5842), .b(net_9695), .c(n5841), .d(net_135) );
na02f01  g2519 ( .o(n8007), .a(n5847), .b(net_9992) );
ao22f01  g2520 ( .o(n8008), .a(n5850), .b(net_9794), .c(n5849_1), .d(net_9893) );
na03f01  g2521 ( .o(n1097), .a(n8008), .b(n8007), .c(n8006_1) );
ao12f01  g2522 ( .o(n8010), .a(n5658), .b(n6160_1), .c(x4694) );
oa12f01  g2523 ( .o(n1102), .a(n8010), .b(n6159), .c(n7772) );
na02f01  g2524 ( .o(n8012), .a(n7937), .b(net_260) );
na02f01  g2525 ( .o(n8013), .a(n7936), .b(net_9790) );
ao22f01  g2526 ( .o(n8014), .a(n7943), .b(_net_10229), .c(n7942), .d(x4041) );
na04f01  g2527 ( .o(n1111), .a(n8014), .b(n8013), .c(n8012), .d(n7939) );
in01f01  g2528 ( .o(n1521), .a(_net_9177) );
in01f01  g2529 ( .o(n8017), .a(_net_9178) );
no02f01  g2530 ( .o(n8018), .a(n8017), .b(n1521) );
in01f01  g2531 ( .o(n8019), .a(n8018) );
na02f01  g2532 ( .o(n8020), .a(n8019), .b(net_9179) );
in01f01  g2533 ( .o(n8021_1), .a(net_9179) );
na02f01  g2534 ( .o(n8022), .a(n8018), .b(n8021_1) );
na02f01  g2535 ( .o(n1116), .a(n8022), .b(n8020) );
in01f01  g2536 ( .o(n8024), .a(net_9182) );
in01f01  g2537 ( .o(n8025), .a(net_9181) );
no02f01  g2538 ( .o(n8026_1), .a(n8025), .b(n8024) );
in01f01  g2539 ( .o(n8027), .a(n8026_1) );
in01f01  g2540 ( .o(n8028), .a(net_9180) );
no02f01  g2541 ( .o(n8029), .a(n8019), .b(n8021_1) );
in01f01  g2542 ( .o(n8030), .a(n8029) );
no02f01  g2543 ( .o(n8031_1), .a(n8030), .b(n8028) );
in01f01  g2544 ( .o(n8032), .a(n8031_1) );
oa12f01  g2545 ( .o(n8033), .a(_net_9183), .b(n8032), .c(n8027) );
in01f01  g2546 ( .o(n8034), .a(_net_9183) );
na03f01  g2547 ( .o(n8035), .a(n8031_1), .b(n8026_1), .c(n8034) );
na02f01  g2548 ( .o(n1125), .a(n8035), .b(n8033) );
oa22f01  g2549 ( .o(n1130), .a(n7367), .b(n6729), .c(n7365_1), .d(n5540) );
ao12f01  g2550 ( .o(n8038), .a(n5658), .b(n7844), .c(_net_259) );
ao22f01  g2551 ( .o(n8039), .a(n7847), .b(x4117), .c(n7846), .d(net_9821) );
na02f01  g2552 ( .o(n1135), .a(n8039), .b(n8038) );
ao22f01  g2553 ( .o(n8041_1), .a(n6599_1), .b(_net_9828), .c(n6572), .d(net_10402) );
no03f01  g2554 ( .o(n8042), .a(n6559), .b(n5549), .c(n5655) );
ao22f01  g2555 ( .o(n8043), .a(n8042), .b(net_10523), .c(n6580), .d(net_9796) );
in01f01  g2556 ( .o(n8044), .a(net_227) );
no03f01  g2557 ( .o(n8045), .a(n6571_1), .b(n6559), .c(x6496) );
in01f01  g2558 ( .o(n8046_1), .a(n8045) );
no02f01  g2559 ( .o(n8047), .a(n6559), .b(n5660) );
ao22f01  g2560 ( .o(n8048), .a(n8047), .b(_net_10062), .c(n6562), .d(_net_200) );
oa12f01  g2561 ( .o(n8049), .a(n8048), .b(n8046_1), .c(n8044) );
na02f01  g2562 ( .o(n8050), .a(n6602), .b(net_9994) );
no03f01  g2563 ( .o(n8051_1), .a(n6559), .b(n5686), .c(x6496) );
ao22f01  g2564 ( .o(n8052), .a(n8051_1), .b(net_90), .c(n6564), .d(net_10075) );
na02f01  g2565 ( .o(n8053), .a(n8052), .b(n8050) );
no02f01  g2566 ( .o(n8054), .a(n8053), .b(n8049) );
ao22f01  g2567 ( .o(n8055_1), .a(n6585), .b(net_9697), .c(n6573), .d(net_9863) );
ao22f01  g2568 ( .o(n8056), .a(n6605), .b(net_10297), .c(n6592), .d(net_10192) );
na02f01  g2569 ( .o(n8057), .a(n8056), .b(n8055_1) );
ao22f01  g2570 ( .o(n8058), .a(n6606), .b(_net_9927), .c(n6555), .d(net_9962) );
ao22f01  g2571 ( .o(n8059_1), .a(n6603), .b(net_10507), .c(n6577), .d(net_9665) );
ao22f01  g2572 ( .o(n8060), .a(n6590), .b(_net_10026), .c(n6584_1), .d(net_9764) );
ao22f01  g2573 ( .o(n8061), .a(n6597), .b(_net_9729), .c(n6582), .d(net_9895) );
na04f01  g2574 ( .o(n8062), .a(n8061), .b(n8060), .c(n8059_1), .d(n8058) );
no02f01  g2575 ( .o(n8063_1), .a(n8062), .b(n8057) );
na04f01  g2576 ( .o(n1140), .a(n8063_1), .b(n8054), .c(n8043), .d(n8041_1) );
na02f01  g2577 ( .o(n8065), .a(n7450), .b(n7398_1) );
in01f01  g2578 ( .o(n8066), .a(n7400) );
na02f01  g2579 ( .o(n8067_1), .a(n7399), .b(n7398_1) );
na03f01  g2580 ( .o(n8068), .a(n8067_1), .b(n7431), .c(n8066) );
na02f01  g2581 ( .o(n8069), .a(n7453), .b(_net_10467) );
na03f01  g2582 ( .o(n1145), .a(n8069), .b(n8068), .c(n8065) );
in01f01  g2583 ( .o(n8071), .a(_net_10417) );
ao12f01  g2584 ( .o(n8072_1), .a(n5658), .b(n6052_1), .c(x5647) );
oa12f01  g2585 ( .o(n1150), .a(n8072_1), .b(n6048), .c(n8071) );
no02f01  g2586 ( .o(n8074), .a(n5498), .b(n5658) );
in01f01  g2587 ( .o(n8075), .a(n8074) );
no02f01  g2588 ( .o(n8076_1), .a(n5495_1), .b(n5658) );
in01f01  g2589 ( .o(n8077), .a(n8076_1) );
no04f01  g2590 ( .o(n8078), .a(n8077), .b(n5501), .c(n5500_1), .d(n5499) );
no03f01  g2591 ( .o(n8079), .a(n5501), .b(x3867), .c(x6157) );
no02f01  g2592 ( .o(n8080), .a(n8079), .b(n5661_1) );
na02f01  g2593 ( .o(n8081_1), .a(n8080), .b(n5504_1) );
no02f01  g2594 ( .o(n8082), .a(n8081_1), .b(n8077) );
ao12f01  g2595 ( .o(n8083), .a(n8078), .b(n8082), .c(net_10530) );
oa12f01  g2596 ( .o(n1155), .a(n8083), .b(n8075), .c(n5626) );
in01f01  g2597 ( .o(n8085), .a(_net_9215) );
in01f01  g2598 ( .o(n8086_1), .a(net_9216) );
in01f01  g2599 ( .o(n8087), .a(_net_9217) );
na03f01  g2600 ( .o(n8088), .a(n8087), .b(n8086_1), .c(n8085) );
in01f01  g2601 ( .o(n8089), .a(_net_9214) );
in01f01  g2602 ( .o(n8090), .a(net_9212) );
in01f01  g2603 ( .o(n8091_1), .a(_net_9211) );
na02f01  g2604 ( .o(n8092), .a(n8091_1), .b(n8090) );
oa12f01  g2605 ( .o(n8093), .a(_net_9213), .b(n8092), .c(net_9210) );
na04f01  g2606 ( .o(n8094), .a(n8093), .b(n8087), .c(n8089), .d(n8086_1) );
na02f01  g2607 ( .o(n8095), .a(n8094), .b(n8088) );
no02f01  g2608 ( .o(n1160), .a(n8095), .b(n6686) );
na02f01  g2609 ( .o(n8097), .a(n7937), .b(net_237) );
na02f01  g2610 ( .o(n8098), .a(n7936), .b(net_9767) );
ao22f01  g2611 ( .o(n8099), .a(n7943), .b(_net_10206), .c(n7942), .d(x5722) );
na04f01  g2612 ( .o(n1165), .a(n8099), .b(n8098), .c(n8097), .d(n7939) );
na02f01  g2613 ( .o(n8101_1), .a(n6147), .b(n6766) );
ao12f01  g2614 ( .o(n8102), .a(n6131_1), .b(n6148), .c(net_9367) );
oa12f01  g2615 ( .o(n1170), .a(n8102), .b(n8101_1), .c(n7088) );
in01f01  g2616 ( .o(n8104), .a(_net_9385) );
in01f01  g2617 ( .o(n8105), .a(_net_9382) );
na02f01  g2618 ( .o(n8106_1), .a(n7446), .b(_net_9381) );
ao12f01  g2619 ( .o(n8107), .a(n8105), .b(n8106_1), .c(n6130) );
ao12f01  g2620 ( .o(n8108), .a(n8107), .b(n8105), .c(n8104) );
in01f01  g2621 ( .o(n8109), .a(n6764) );
in01f01  g2622 ( .o(n8110), .a(x589) );
no03f01  g2623 ( .o(n8111_1), .a(n8110), .b(_net_9164), .c(x3653) );
no04f01  g2624 ( .o(n8112), .a(n8111_1), .b(n8109), .c(net_9163), .d(net_9289) );
ao12f01  g2625 ( .o(n1179), .a(n5658), .b(n8112), .c(n8108) );
in01f01  g2626 ( .o(n8114), .a(net_9509) );
no03f01  g2627 ( .o(n8115), .a(_net_8955), .b(_net_9062), .c(n5738) );
na02f01  g2628 ( .o(n8116_1), .a(n8115), .b(n5697) );
no02f01  g2629 ( .o(n8117), .a(n8115), .b(_net_9421) );
no02f01  g2630 ( .o(n8118), .a(n8117), .b(n5697) );
ao22f01  g2631 ( .o(n8119), .a(n8118), .b(x2968), .c(n8117), .d(_net_9394) );
oa12f01  g2632 ( .o(n1183), .a(n8119), .b(n8116_1), .c(n8114) );
in01f01  g2633 ( .o(n8121), .a(_net_10411) );
ao12f01  g2634 ( .o(n8122), .a(n5658), .b(n6052_1), .c(x6028) );
oa12f01  g2635 ( .o(n1188), .a(n8122), .b(n6048), .c(n8121) );
no04f01  g2636 ( .o(n1193), .a(net_9273), .b(net_9274), .c(_net_9272), .d(n5658) );
oa22f01  g2637 ( .o(n8125_1), .a(n7778_1), .b(n6723_1), .c(n7769), .d(n6720) );
no02f01  g2638 ( .o(n8126), .a(_net_10154), .b(_net_9730) );
no02f01  g2639 ( .o(n8127), .a(n7785), .b(n6729) );
no02f01  g2640 ( .o(n8128), .a(n7782_1), .b(n6727) );
no02f01  g2641 ( .o(n8129), .a(_net_10153), .b(_net_9729) );
in01f01  g2642 ( .o(n8130_1), .a(n8129) );
ao12f01  g2643 ( .o(n8131), .a(n8127), .b(n8130_1), .c(n8128) );
no02f01  g2644 ( .o(n8132), .a(n8131), .b(n8126) );
oa22f01  g2645 ( .o(n8133), .a(n8132), .b(n8125_1), .c(_net_10155), .d(_net_9731) );
no02f01  g2646 ( .o(n8134), .a(n6736), .b(n7767) );
no02f01  g2647 ( .o(n8135_1), .a(_net_9732), .b(_net_10156) );
no02f01  g2648 ( .o(n8136), .a(n8135_1), .b(n8134) );
in01f01  g2649 ( .o(n8137), .a(n8136) );
ao12f01  g2650 ( .o(n8138), .a(n6746), .b(n8137), .c(n8133) );
oa12f01  g2651 ( .o(n8139), .a(n8138), .b(n8137), .c(n8133) );
no02f01  g2652 ( .o(n8140_1), .a(_net_10152), .b(_net_10153) );
in01f01  g2653 ( .o(n8141), .a(n8140_1) );
no02f01  g2654 ( .o(n8142), .a(n8141), .b(_net_10154) );
na02f01  g2655 ( .o(n8143), .a(n8142), .b(n7769) );
no02f01  g2656 ( .o(n8144), .a(n8143), .b(_net_10156) );
in01f01  g2657 ( .o(n8145_1), .a(n8144) );
na02f01  g2658 ( .o(n8146), .a(n8143), .b(_net_10156) );
na02f01  g2659 ( .o(n8147), .a(n8146), .b(n8145_1) );
ao22f01  g2660 ( .o(n8148), .a(n8147), .b(n6750), .c(n6760), .d(_net_10156) );
na02f01  g2661 ( .o(n1198), .a(n8148), .b(n8139) );
ao12f01  g2662 ( .o(n8150_1), .a(n5658), .b(n6875_1), .c(net_251) );
ao22f01  g2663 ( .o(n8151), .a(n6878), .b(x4781), .c(n6877), .d(net_9912) );
na02f01  g2664 ( .o(n1203), .a(n8151), .b(n8150_1) );
in01f01  g2665 ( .o(n8153), .a(net_9948) );
oa22f01  g2666 ( .o(n1208), .a(n5694), .b(n8153), .c(n5692), .d(n5567_1) );
no02f01  g2667 ( .o(n8155_1), .a(_net_9931), .b(_net_10367) );
in01f01  g2668 ( .o(n8156), .a(n8155_1) );
no02f01  g2669 ( .o(n8157), .a(n5722), .b(n7010) );
no02f01  g2670 ( .o(n8158), .a(n7012_1), .b(n5721) );
ao12f01  g2671 ( .o(n8159), .a(n8157), .b(n8158), .c(n8156) );
in01f01  g2672 ( .o(n8160_1), .a(n8159) );
no02f01  g2673 ( .o(n8161), .a(_net_10366), .b(_net_9930) );
no02f01  g2674 ( .o(n8162), .a(n7024), .b(n5711) );
in01f01  g2675 ( .o(n8163), .a(n8162) );
no02f01  g2676 ( .o(n8164), .a(n7015), .b(n5710_1) );
in01f01  g2677 ( .o(n8165_1), .a(n8164) );
na02f01  g2678 ( .o(n8166), .a(n8165_1), .b(n8163) );
no02f01  g2679 ( .o(n8167), .a(_net_10364), .b(_net_9928) );
no02f01  g2680 ( .o(n8168), .a(n7031), .b(n5706) );
no02f01  g2681 ( .o(n8169), .a(n5707), .b(n7029) );
no02f01  g2682 ( .o(n8170_1), .a(_net_10363), .b(_net_9927) );
in01f01  g2683 ( .o(n8171), .a(n8170_1) );
ao12f01  g2684 ( .o(n8172), .a(n8168), .b(n8171), .c(n8169) );
no02f01  g2685 ( .o(n8173), .a(n8172), .b(n8167) );
oa22f01  g2686 ( .o(n8174), .a(n8173), .b(n8166), .c(_net_10365), .d(_net_9929) );
no02f01  g2687 ( .o(n8175_1), .a(n8174), .b(n8161) );
ao12f01  g2688 ( .o(n8176), .a(n8160_1), .b(n8175_1), .c(n8156) );
in01f01  g2689 ( .o(n8177), .a(n8176) );
no02f01  g2690 ( .o(n8178), .a(n5718), .b(n7007_1) );
no02f01  g2691 ( .o(n8179), .a(_net_9932), .b(_net_10368) );
no02f01  g2692 ( .o(n8180_1), .a(n8179), .b(n8178) );
in01f01  g2693 ( .o(n8181), .a(_net_9938) );
oa12f01  g2694 ( .o(n8182), .a(net_10385), .b(n6165), .c(_net_8830) );
no03f01  g2695 ( .o(n8183), .a(n8182), .b(n8181), .c(net_10409) );
in01f01  g2696 ( .o(n8184), .a(n8183) );
ao12f01  g2697 ( .o(n8185_1), .a(n8184), .b(n8180_1), .c(n8177) );
oa12f01  g2698 ( .o(n8186), .a(n8185_1), .b(n8180_1), .c(n8177) );
no02f01  g2699 ( .o(n8187), .a(_net_10362), .b(_net_10363) );
in01f01  g2700 ( .o(n8188), .a(n8187) );
no02f01  g2701 ( .o(n8189), .a(n8188), .b(_net_10364) );
na02f01  g2702 ( .o(n8190_1), .a(n8189), .b(n7015) );
no02f01  g2703 ( .o(n8191), .a(n8190_1), .b(_net_10366) );
in01f01  g2704 ( .o(n8192), .a(n8191) );
no02f01  g2705 ( .o(n8193), .a(n8192), .b(_net_10367) );
in01f01  g2706 ( .o(n8194), .a(n8193) );
no02f01  g2707 ( .o(n8195_1), .a(n8194), .b(_net_10368) );
in01f01  g2708 ( .o(n8196), .a(n8195_1) );
na02f01  g2709 ( .o(n8197), .a(n8194), .b(_net_10368) );
na02f01  g2710 ( .o(n8198), .a(n8197), .b(n8196) );
in01f01  g2711 ( .o(n8199), .a(net_10409) );
no02f01  g2712 ( .o(n8200_1), .a(n8181), .b(n8199) );
in01f01  g2713 ( .o(n8201), .a(n8182) );
no03f01  g2714 ( .o(n8202), .a(n8201), .b(n8181), .c(net_10409) );
ao22f01  g2715 ( .o(n8203), .a(n8202), .b(_net_10368), .c(n8200_1), .d(n8198) );
na02f01  g2716 ( .o(n1213), .a(n8203), .b(n8186) );
na02f01  g2717 ( .o(n8205_1), .a(n6056), .b(net_237) );
na02f01  g2718 ( .o(n8206), .a(n6055), .b(net_9965) );
ao22f01  g2719 ( .o(n8207), .a(n6062_1), .b(x5722), .c(n6060), .d(_net_10416) );
na04f01  g2720 ( .o(n1222), .a(n8207), .b(n8206), .c(n8205_1), .d(n6058) );
in01f01  g2721 ( .o(n8209), .a(_net_10434) );
no02f01  g2722 ( .o(n8210_1), .a(_net_10472), .b(n8209) );
no02f01  g2723 ( .o(n8211), .a(n7413_1), .b(_net_10434) );
in01f01  g2724 ( .o(n8212), .a(n8211) );
in01f01  g2725 ( .o(n8213), .a(_net_10433) );
no02f01  g2726 ( .o(n8214_1), .a(n8213), .b(_net_10471) );
ao12f01  g2727 ( .o(n8215), .a(n8210_1), .b(n8214_1), .c(n8212) );
no02f01  g2728 ( .o(n8216), .a(_net_10433), .b(n7415) );
in01f01  g2729 ( .o(n8217), .a(n8216) );
no02f01  g2730 ( .o(n8218), .a(_net_10432), .b(n7433) );
in01f01  g2731 ( .o(n8219_1), .a(_net_10432) );
no02f01  g2732 ( .o(n8220), .a(_net_10469), .b(n7361) );
in01f01  g2733 ( .o(n8221), .a(n8220) );
oa12f01  g2734 ( .o(n8222), .a(n8219_1), .b(n8221), .c(_net_10470) );
oa12f01  g2735 ( .o(n8223_1), .a(_net_10470), .b(n8221), .c(n8219_1) );
na02f01  g2736 ( .o(n8224), .a(n8223_1), .b(n8222) );
no02f01  g2737 ( .o(n8225), .a(n7388), .b(_net_10431) );
in01f01  g2738 ( .o(n8226), .a(n8225) );
in01f01  g2739 ( .o(n8227_1), .a(_net_10430) );
no02f01  g2740 ( .o(n8228), .a(n8227_1), .b(_net_10468) );
no02f01  g2741 ( .o(n8229), .a(n7398_1), .b(_net_10429) );
no02f01  g2742 ( .o(n8230), .a(_net_10430), .b(n7395) );
no02f01  g2743 ( .o(n8231_1), .a(n8230), .b(n8229) );
no02f01  g2744 ( .o(n8232), .a(n8231_1), .b(n8228) );
in01f01  g2745 ( .o(n8233), .a(n8232) );
na02f01  g2746 ( .o(n8234), .a(n8233), .b(n8226) );
oa12f01  g2747 ( .o(n8235_1), .a(n8224), .b(n8234), .c(n8218) );
na02f01  g2748 ( .o(n8236), .a(n8235_1), .b(n8217) );
no02f01  g2749 ( .o(n8237), .a(n8236), .b(n8211) );
in01f01  g2750 ( .o(n8238), .a(n8237) );
no02f01  g2751 ( .o(n8239), .a(n7380), .b(_net_10435) );
in01f01  g2752 ( .o(n8240_1), .a(_net_10435) );
no02f01  g2753 ( .o(n8241), .a(_net_10473), .b(n8240_1) );
no02f01  g2754 ( .o(n8242), .a(n8241), .b(n8239) );
na03f01  g2755 ( .o(n8243), .a(n8242), .b(n8238), .c(n8215) );
in01f01  g2756 ( .o(n8244), .a(n8215) );
in01f01  g2757 ( .o(n8245_1), .a(n8242) );
oa12f01  g2758 ( .o(n8246), .a(n8245_1), .b(n8237), .c(n8244) );
na02f01  g2759 ( .o(n1227), .a(n8246), .b(n8243) );
in01f01  g2760 ( .o(n8248), .a(_net_9751) );
oa22f01  g2761 ( .o(n1232), .a(n7367), .b(n8248), .c(n7365_1), .d(n5609) );
ao22f01  g2762 ( .o(n8250_1), .a(n5842), .b(net_9757), .c(n5841), .d(_net_8833) );
na02f01  g2763 ( .o(n8251), .a(n5847), .b(_net_10054) );
ao22f01  g2764 ( .o(n8252), .a(n5850), .b(net_9856), .c(n5849_1), .d(net_9955) );
na03f01  g2765 ( .o(n1242), .a(n8252), .b(n8251), .c(n8250_1) );
in01f01  g2766 ( .o(n8254), .a(net_206) );
in01f01  g2767 ( .o(n8255_1), .a(net_205) );
in01f01  g2768 ( .o(n8256), .a(net_204) );
in01f01  g2769 ( .o(n8257), .a(net_203) );
in01f01  g2770 ( .o(n8258), .a(_net_202) );
in01f01  g2771 ( .o(n8259), .a(_net_201) );
in01f01  g2772 ( .o(n8260_1), .a(_net_200) );
in01f01  g2773 ( .o(n8261), .a(_net_199) );
na02f01  g2774 ( .o(n8262), .a(_net_198), .b(net_197) );
no02f01  g2775 ( .o(n8263), .a(n8262), .b(n8261) );
in01f01  g2776 ( .o(n8264_1), .a(n8263) );
no02f01  g2777 ( .o(n8265), .a(n8264_1), .b(n8260_1) );
in01f01  g2778 ( .o(n8266), .a(n8265) );
no02f01  g2779 ( .o(n8267), .a(n8266), .b(n8259) );
in01f01  g2780 ( .o(n8268_1), .a(n8267) );
no02f01  g2781 ( .o(n8269), .a(n8268_1), .b(n8258) );
in01f01  g2782 ( .o(n8270), .a(n8269) );
no02f01  g2783 ( .o(n8271), .a(n8270), .b(n8257) );
in01f01  g2784 ( .o(n8272_1), .a(n8271) );
no02f01  g2785 ( .o(n8273), .a(n8272_1), .b(n8256) );
in01f01  g2786 ( .o(n8274), .a(n8273) );
no02f01  g2787 ( .o(n8275), .a(n8274), .b(n8255_1) );
na02f01  g2788 ( .o(n8276_1), .a(n8275), .b(net_206) );
in01f01  g2789 ( .o(n8277), .a(n8276_1) );
oa12f01  g2790 ( .o(n8278), .a(n573), .b(n8275), .c(net_206) );
in01f01  g2791 ( .o(n8279), .a(_net_9268) );
na02f01  g2792 ( .o(n8280), .a(n8279), .b(n5914) );
oa22f01  g2793 ( .o(n1247), .a(n8280), .b(n8254), .c(n8278), .d(n8277) );
in01f01  g2794 ( .o(n8282), .a(net_10084) );
oa22f01  g2795 ( .o(n1252), .a(n6989_1), .b(n5546), .c(n6988), .d(n8282) );
in01f01  g2796 ( .o(n8284), .a(net_213) );
ao22f01  g2797 ( .o(n8285), .a(n8047), .b(net_10063), .c(n6564), .d(net_10085) );
oa12f01  g2798 ( .o(n8286_1), .a(n8285), .b(n6563), .c(n8284) );
ao22f01  g2799 ( .o(n8287), .a(n6592), .b(net_10186), .c(n6580), .d(net_9813) );
ao22f01  g2800 ( .o(n8288), .a(n6577), .b(net_9682), .c(n6572), .d(net_10396) );
na02f01  g2801 ( .o(n8289), .a(n8288), .b(n8287) );
no02f01  g2802 ( .o(n8290), .a(n8289), .b(n8286_1) );
ao22f01  g2803 ( .o(n8291_1), .a(n6606), .b(_net_9943), .c(n6597), .d(_net_9745) );
ao22f01  g2804 ( .o(n8292), .a(n6585), .b(net_9714), .c(n6584_1), .d(net_9781) );
na02f01  g2805 ( .o(n8293), .a(n6555), .b(net_9979) );
na02f01  g2806 ( .o(n8294), .a(n6602), .b(net_10011) );
na02f01  g2807 ( .o(n8295), .a(n8294), .b(n8293) );
na02f01  g2808 ( .o(n8296_1), .a(n6573), .b(net_9880) );
oa12f01  g2809 ( .o(n8297), .a(n8296_1), .b(n6591), .c(n5829) );
in01f01  g2810 ( .o(n8298), .a(net_10501) );
in01f01  g2811 ( .o(n8299), .a(n6603) );
oa22f01  g2812 ( .o(n8300), .a(n8299), .b(n8298), .c(n6600), .d(n5799) );
in01f01  g2813 ( .o(n8301_1), .a(net_10291) );
in01f01  g2814 ( .o(n8302), .a(n6605) );
na02f01  g2815 ( .o(n8303), .a(n6582), .b(net_9912) );
oa12f01  g2816 ( .o(n8304), .a(n8303), .b(n8302), .c(n8301_1) );
no04f01  g2817 ( .o(n8305_1), .a(n8304), .b(n8300), .c(n8297), .d(n8295) );
na04f01  g2818 ( .o(n1257), .a(n8305_1), .b(n8292), .c(n8291_1), .d(n8290) );
in01f01  g2819 ( .o(n8307), .a(_net_10319) );
ao12f01  g2820 ( .o(n8308), .a(n5658), .b(n5774), .c(x5225) );
oa12f01  g2821 ( .o(n1262), .a(n8308), .b(n5770), .c(n8307) );
in01f01  g2822 ( .o(n8310_1), .a(net_10181) );
oa22f01  g2823 ( .o(n1267), .a(n7956), .b(n5525), .c(n7955), .d(n8310_1) );
ao12f01  g2824 ( .o(n8312), .a(n5658), .b(n6532), .c(_net_261) );
ao22f01  g2825 ( .o(n8313), .a(n6535), .b(x3949), .c(n6534), .d(net_10021) );
na02f01  g2826 ( .o(n1272), .a(n8313), .b(n8312) );
ao22f01  g2827 ( .o(n8315_1), .a(n5842), .b(net_9723), .c(n5841), .d(_net_163) );
na02f01  g2828 ( .o(n8316), .a(n5847), .b(net_10020) );
ao22f01  g2829 ( .o(n8317), .a(n5850), .b(net_9822), .c(n5849_1), .d(net_9921) );
na03f01  g2830 ( .o(n1277), .a(n8317), .b(n8316), .c(n8315_1) );
na02f01  g2831 ( .o(n8319), .a(net_10291), .b(net_10299) );
ao22f01  g2832 ( .o(n8320_1), .a(net_10292), .b(net_10300), .c(net_10298), .d(net_10290) );
ao22f01  g2833 ( .o(n8321), .a(net_10287), .b(net_10294), .c(net_10297), .d(net_10290) );
ao22f01  g2834 ( .o(n8322), .a(net_10288), .b(net_10295), .c(net_10289), .d(net_10296) );
na04f01  g2835 ( .o(n1286), .a(n8322), .b(n8321), .c(n8320_1), .d(n8319) );
no02f01  g2836 ( .o(n8324), .a(n8230), .b(n8228) );
na02f01  g2837 ( .o(n8325_1), .a(n8324), .b(n8229) );
in01f01  g2838 ( .o(n8326), .a(n8229) );
oa12f01  g2839 ( .o(n8327), .a(n8326), .b(n8230), .c(n8228) );
na02f01  g2840 ( .o(n1291), .a(n8327), .b(n8325_1) );
in01f01  g2841 ( .o(n8329), .a(net_9760) );
in01f01  g2842 ( .o(n8330_1), .a(net_9759) );
na02f01  g2843 ( .o(n1301), .a(n8330_1), .b(n8329) );
in01f01  g2844 ( .o(n8332), .a(_net_9320) );
in01f01  g2845 ( .o(n8333), .a(_net_9312) );
in01f01  g2846 ( .o(n8334), .a(_net_9326) );
no02f01  g2847 ( .o(n8335_1), .a(n8334), .b(n8333) );
no02f01  g2848 ( .o(n8336), .a(_net_9326), .b(_net_9312) );
no02f01  g2849 ( .o(n8337), .a(n8336), .b(n8335_1) );
no02f01  g2850 ( .o(n8338), .a(n8337), .b(net_9152) );
in01f01  g2851 ( .o(n8339_1), .a(net_9152) );
no03f01  g2852 ( .o(n8340), .a(n8336), .b(n8335_1), .c(n8339_1) );
no02f01  g2853 ( .o(n8341), .a(n8340), .b(n8338) );
ao12f01  g2854 ( .o(n8342), .a(n7883), .b(n8341), .c(n7923) );
oa12f01  g2855 ( .o(n1306), .a(n8342), .b(n7925_1), .c(n8332) );
in01f01  g2856 ( .o(n8344_1), .a(_net_9191) );
in01f01  g2857 ( .o(n8345), .a(_net_9185) );
no02f01  g2858 ( .o(n8346), .a(n7698), .b(_net_9167) );
na03f01  g2859 ( .o(n8347), .a(n8346), .b(n7702), .c(n8345) );
in01f01  g2860 ( .o(n8348), .a(n8346) );
na03f01  g2861 ( .o(n8349_1), .a(n8348), .b(n7702), .c(n8345) );
oa22f01  g2862 ( .o(n1315), .a(n8349_1), .b(n8024), .c(n8347), .d(n8344_1) );
oa22f01  g2863 ( .o(n1320), .a(n5694), .b(n5718), .c(n5692), .d(n5606) );
ao12f01  g2864 ( .o(n8352), .a(n5658), .b(n6875_1), .c(net_241) );
ao22f01  g2865 ( .o(n8353), .a(n6878), .b(x5498), .c(n6877), .d(net_9902) );
na02f01  g2866 ( .o(n1325), .a(n8353), .b(n8352) );
na02f01  g2867 ( .o(n8355), .a(n6038), .b(_net_231) );
na02f01  g2868 ( .o(n8356), .a(n6037_1), .b(net_9860) );
ao22f01  g2869 ( .o(n8357), .a(n6044), .b(x6102), .c(n6042_1), .d(_net_10305) );
na04f01  g2870 ( .o(n1330), .a(n8357), .b(n8356), .c(n8355), .d(n6040) );
na02f01  g2871 ( .o(n8359), .a(n6056), .b(net_250) );
na02f01  g2872 ( .o(n8360), .a(n6055), .b(net_9978) );
ao22f01  g2873 ( .o(n8361), .a(n6062_1), .b(x4851), .c(n6060), .d(_net_10429) );
na04f01  g2874 ( .o(n1339), .a(n8361), .b(n8360), .c(n8359), .d(n6058) );
in01f01  g2875 ( .o(n8363_1), .a(net_9924) );
oa22f01  g2876 ( .o(n1344), .a(n5694), .b(n8363_1), .c(n5692), .d(n5570) );
ao22f01  g2877 ( .o(n8365), .a(n5842), .b(net_9715), .c(n5841), .d(_net_155) );
na02f01  g2878 ( .o(n8366), .a(n5847), .b(net_10012) );
ao22f01  g2879 ( .o(n8367), .a(n5850), .b(net_9814), .c(n5849_1), .d(net_9913) );
na03f01  g2880 ( .o(n1349), .a(n8367), .b(n8366), .c(n8365) );
in01f01  g2881 ( .o(n8369), .a(net_9670) );
in01f01  g2882 ( .o(n8370), .a(n6577) );
ao22f01  g2883 ( .o(n8371), .a(n6564), .b(net_10080), .c(n6562), .d(net_205) );
oa12f01  g2884 ( .o(n8372_1), .a(n8371), .b(n8370), .c(n8369) );
ao22f01  g2885 ( .o(n8373), .a(n6597), .b(_net_9734), .c(n6584_1), .d(net_9769) );
na02f01  g2886 ( .o(n8374), .a(n6582), .b(net_9900) );
na02f01  g2887 ( .o(n8375), .a(n6602), .b(net_9999) );
na03f01  g2888 ( .o(n8376_1), .a(n8375), .b(n8374), .c(n8373) );
no02f01  g2889 ( .o(n8377), .a(n8376_1), .b(n8372_1) );
na02f01  g2890 ( .o(n8378), .a(n6555), .b(net_9967) );
na02f01  g2891 ( .o(n8379), .a(n6573), .b(net_9868) );
na02f01  g2892 ( .o(n8380_1), .a(n8379), .b(n8378) );
ao12f01  g2893 ( .o(n8381), .a(n8380_1), .b(n6590), .c(_net_10031) );
ao22f01  g2894 ( .o(n8382), .a(n6606), .b(_net_9932), .c(n6580), .d(net_9801) );
ao22f01  g2895 ( .o(n8383), .a(n6599_1), .b(_net_9833), .c(n6585), .d(net_9702) );
na04f01  g2896 ( .o(n1354), .a(n8383), .b(n8382), .c(n8381), .d(n8377) );
na02f01  g2897 ( .o(n8385), .a(n7353), .b(x5143) );
na02f01  g2898 ( .o(n8386), .a(n7352), .b(net_9677) );
ao22f01  g2899 ( .o(n8387), .a(n7358), .b(net_246), .c(n7357), .d(_net_10110) );
na04f01  g2900 ( .o(n1359), .a(n8387), .b(n8386), .c(n8385), .d(n7355_1) );
in01f01  g2901 ( .o(n8389_1), .a(_net_9186) );
oa22f01  g2902 ( .o(n1369), .a(n8349_1), .b(n1521), .c(n8347), .d(n8389_1) );
ao22f01  g2903 ( .o(n8391), .a(n5842), .b(net_9718), .c(n5841), .d(_net_158) );
na02f01  g2904 ( .o(n8392), .a(n5847), .b(net_10015) );
ao22f01  g2905 ( .o(n8393), .a(n5850), .b(net_9817), .c(n5849_1), .d(net_9916) );
na03f01  g2906 ( .o(n1374), .a(n8393), .b(n8392), .c(n8391) );
in01f01  g2907 ( .o(n8395), .a(_net_10336) );
ao12f01  g2908 ( .o(n8396), .a(n5658), .b(n5774), .c(x3889) );
oa12f01  g2909 ( .o(n1379), .a(n8396), .b(n5770), .c(n8395) );
na03f01  g2910 ( .o(n8398), .a(n5880), .b(n5879), .c(_net_9536) );
in01f01  g2911 ( .o(n8399_1), .a(_net_9250) );
na02f01  g2912 ( .o(n8400), .a(n5887), .b(n8399_1) );
in01f01  g2913 ( .o(n8401), .a(n8400) );
no02f01  g2914 ( .o(n8402), .a(net_9542), .b(n7979) );
na02f01  g2915 ( .o(n8403), .a(n5489), .b(_net_9536) );
na02f01  g2916 ( .o(n8404_1), .a(n5890), .b(n8399_1) );
in01f01  g2917 ( .o(n8405), .a(_net_9503) );
na02f01  g2918 ( .o(n8406), .a(n8405), .b(_net_9536) );
oa22f01  g2919 ( .o(n8407), .a(n8406), .b(n8404_1), .c(n8403), .d(n5871) );
ao12f01  g2920 ( .o(n8408), .a(n8407), .b(n8402), .c(n8401) );
in01f01  g2921 ( .o(n8409_1), .a(n5856) );
oa12f01  g2922 ( .o(n8410), .a(n8409_1), .b(n5854), .c(n7979) );
oa12f01  g2923 ( .o(n8411), .a(x6599), .b(_net_9537), .c(_net_9536) );
na02f01  g2924 ( .o(n8412), .a(n8411), .b(n5866) );
no02f01  g2925 ( .o(n8413), .a(n8403), .b(_net_9250) );
ao22f01  g2926 ( .o(n8414_1), .a(n8413), .b(n8412), .c(n8410), .d(n5859) );
na03f01  g2927 ( .o(n1384), .a(n8414_1), .b(n8408), .c(n8398) );
in01f01  g2928 ( .o(n8416), .a(net_228) );
na03f01  g2929 ( .o(n8417), .a(n8045), .b(n5663), .c(x6599) );
oa12f01  g2930 ( .o(n8418), .a(x6599), .b(n8046_1), .c(n5664) );
oa22f01  g2931 ( .o(n1392), .a(n8418), .b(n8416), .c(n8417), .d(n5573) );
in01f01  g2932 ( .o(n8420), .a(net_9653) );
na02f01  g2933 ( .o(n8421), .a(net_9654), .b(n6514) );
in01f01  g2934 ( .o(n8422), .a(net_9654) );
na02f01  g2935 ( .o(n8423), .a(n8422), .b(net_313) );
na04f01  g2936 ( .o(n8424_1), .a(n8423), .b(n8421), .c(net_9652), .d(n8420) );
no02f01  g2937 ( .o(n8425), .a(net_9651), .b(net_313) );
in01f01  g2938 ( .o(n8426), .a(net_9651) );
no02f01  g2939 ( .o(n8427), .a(n8426), .b(n6514) );
no02f01  g2940 ( .o(n8428), .a(n8427), .b(n8425) );
no02f01  g2941 ( .o(n8429_1), .a(net_9655), .b(n6514) );
in01f01  g2942 ( .o(n8430), .a(net_9655) );
no02f01  g2943 ( .o(n8431), .a(n8430), .b(net_313) );
no03f01  g2944 ( .o(n8432), .a(net_9657), .b(net_9656), .c(net_9650) );
oa12f01  g2945 ( .o(n8433_1), .a(n8432), .b(n8431), .c(n8429_1) );
no03f01  g2946 ( .o(n1401), .a(n8433_1), .b(n8428), .c(n8424_1) );
no02f01  g2947 ( .o(n8435), .a(n7025), .b(n7019) );
in01f01  g2948 ( .o(n8436), .a(n8435) );
na02f01  g2949 ( .o(n8437), .a(n8436), .b(n7035) );
na02f01  g2950 ( .o(n8438_1), .a(n8435), .b(n7034_1) );
na02f01  g2951 ( .o(n1406), .a(n8438_1), .b(n8437) );
in01f01  g2952 ( .o(n8440), .a(net_10180) );
oa22f01  g2953 ( .o(n1415), .a(n7956), .b(n5615), .c(n7955), .d(n8440) );
in01f01  g2954 ( .o(n8442), .a(_net_10126) );
ao12f01  g2955 ( .o(n8443_1), .a(n5658), .b(n6160_1), .c(x3889) );
oa12f01  g2956 ( .o(n1420), .a(n8443_1), .b(n6159), .c(n8442) );
oa22f01  g2957 ( .o(n1425), .a(n5694), .b(n5721), .c(n5692), .d(n5561) );
in01f01  g2958 ( .o(n8446), .a(_net_9242) );
na02f01  g2959 ( .o(n6033), .a(n8446), .b(n6475) );
na04f01  g2960 ( .o(n8448), .a(n7852), .b(n6520), .c(n6507_1), .d(n6504) );
no02f01  g2961 ( .o(n8449), .a(n8448), .b(n6033) );
no02f01  g2962 ( .o(n8450), .a(_net_9240), .b(_net_9239) );
in01f01  g2963 ( .o(n8451), .a(n8450) );
no02f01  g2964 ( .o(n8452_1), .a(_net_9237), .b(_net_9238) );
na02f01  g2965 ( .o(n8453), .a(n8452_1), .b(n6511) );
no03f01  g2966 ( .o(n8454), .a(n8453), .b(n8451), .c(_net_9241) );
na02f01  g2967 ( .o(n1430), .a(n8454), .b(n8449) );
no02f01  g2968 ( .o(n8456), .a(n7071), .b(_net_9293) );
in01f01  g2969 ( .o(n8457_1), .a(n8456) );
oa12f01  g2970 ( .o(n8458), .a(n8457_1), .b(n7573), .c(_net_9292) );
na02f01  g2971 ( .o(n8459), .a(n7071), .b(_net_9293) );
na02f01  g2972 ( .o(n8460), .a(n5916), .b(_net_9291) );
oa12f01  g2973 ( .o(n8461), .a(n8460), .b(n7593), .c(_net_167) );
oa12f01  g2974 ( .o(n8462_1), .a(n8461), .b(n5916), .c(_net_9291) );
no02f01  g2975 ( .o(n8463), .a(_net_170), .b(n7073_1) );
ao12f01  g2976 ( .o(n8464), .a(n8463), .b(n7573), .c(_net_9292) );
ao22f01  g2977 ( .o(n8465), .a(n8464), .b(n8462_1), .c(n8459), .d(n8458) );
in01f01  g2978 ( .o(n8466), .a(_net_173) );
ao22f01  g2979 ( .o(n8467_1), .a(_net_9297), .b(n7554), .c(n8466), .d(_net_9296) );
in01f01  g2980 ( .o(n8468), .a(_net_171) );
in01f01  g2981 ( .o(n8469), .a(_net_9295) );
no02f01  g2982 ( .o(n8470), .a(n8469), .b(_net_172) );
ao12f01  g2983 ( .o(n8471), .a(n8470), .b(n8468), .c(_net_9294) );
na02f01  g2984 ( .o(n8472_1), .a(n8471), .b(n8467_1) );
ao22f01  g2985 ( .o(n8473), .a(n7552_1), .b(_net_174), .c(_net_173), .d(n7545) );
ao12f01  g2986 ( .o(n8474), .a(n8473), .b(_net_9297), .c(n7554) );
no02f01  g2987 ( .o(n8475), .a(_net_9295), .b(n5975) );
in01f01  g2988 ( .o(n8476), .a(n8475) );
na02f01  g2989 ( .o(n8477_1), .a(_net_171), .b(n7605_1) );
oa12f01  g2990 ( .o(n8478), .a(n8476), .b(n8477_1), .c(n8470) );
ao12f01  g2991 ( .o(n8479), .a(n8474), .b(n8478), .c(n8467_1) );
oa12f01  g2992 ( .o(n8480), .a(n8479), .b(n8472_1), .c(n8465) );
no02f01  g2993 ( .o(n8481), .a(_net_175), .b(n7536) );
no02f01  g2994 ( .o(n8482_1), .a(n7529_1), .b(_net_176) );
no02f01  g2995 ( .o(n8483), .a(_net_177), .b(n7516) );
no03f01  g2996 ( .o(n8484), .a(n8483), .b(n8482_1), .c(n8481) );
in01f01  g2997 ( .o(n8485), .a(n8482_1) );
no02f01  g2998 ( .o(n8486_1), .a(_net_9299), .b(n5990) );
no02f01  g2999 ( .o(n8487), .a(n5989), .b(_net_9298) );
ao12f01  g3000 ( .o(n8488), .a(n8486_1), .b(n8487), .c(n8485) );
no02f01  g3001 ( .o(n8489), .a(n5983_1), .b(_net_9300) );
no02f01  g3002 ( .o(n8490), .a(n8489), .b(_net_182) );
oa12f01  g3003 ( .o(n8491_1), .a(n8490), .b(n8488), .c(n8483) );
ao12f01  g3004 ( .o(n1435), .a(n8491_1), .b(n8484), .c(n8480) );
na02f01  g3005 ( .o(n8493), .a(n7358), .b(_net_234) );
na02f01  g3006 ( .o(n8494), .a(n7352), .b(net_9665) );
ao22f01  g3007 ( .o(n8495), .a(n7357), .b(_net_10098), .c(n7353), .d(x5901) );
na04f01  g3008 ( .o(n1444), .a(n8495), .b(n8494), .c(n8493), .d(n7355_1) );
no03f01  g3009 ( .o(n8497), .a(n6474_1), .b(n6475), .c(n6463) );
na02f01  g3010 ( .o(n8498), .a(n6471), .b(_net_9245) );
ao12f01  g3011 ( .o(n8499), .a(n8498), .b(n7863), .c(n7852) );
na03f01  g3012 ( .o(n8500), .a(n6860), .b(_net_9236), .c(_net_9245) );
oa12f01  g3013 ( .o(n8501_1), .a(n8500), .b(n8498), .c(n7862_1) );
na03f01  g3014 ( .o(n8502), .a(n6850), .b(n6486), .c(_net_9245) );
no03f01  g3015 ( .o(n8503), .a(n6136), .b(n6491), .c(n6475) );
no03f01  g3016 ( .o(n8504), .a(_net_9169), .b(n8446), .c(n6475) );
no03f01  g3017 ( .o(n8505_1), .a(_net_9209), .b(n6520), .c(n6475) );
no03f01  g3018 ( .o(n8506), .a(n8505_1), .b(n8504), .c(n8503) );
no03f01  g3019 ( .o(n8507), .a(n6495), .b(_net_9172), .c(n6475) );
in01f01  g3020 ( .o(n8508), .a(_net_9169) );
in01f01  g3021 ( .o(n8509), .a(_net_9244) );
ao12f01  g3022 ( .o(n8510_1), .a(n8509), .b(n8508), .c(n6475) );
no03f01  g3023 ( .o(n8511), .a(n6489_1), .b(n6475), .c(_net_9171) );
no04f01  g3024 ( .o(n8512), .a(n8511), .b(n8510_1), .c(n8507), .d(n6476) );
na03f01  g3025 ( .o(n8513), .a(n8512), .b(n8506), .c(n8502) );
no04f01  g3026 ( .o(n8514), .a(n8513), .b(n8501_1), .c(n8499), .d(n8497) );
no02f01  g3027 ( .o(n1449), .a(n8514), .b(n6526_1) );
na02f01  g3028 ( .o(n8516), .a(n6020), .b(n7072) );
oa12f01  g3029 ( .o(n1454), .a(n8516), .b(n6020), .c(n7071) );
ao12f01  g3030 ( .o(n8518), .a(n7572), .b(n6028_1), .c(n6625) );
oa12f01  g3031 ( .o(n1459), .a(n8518), .b(n6022), .c(n7573) );
ao12f01  g3032 ( .o(n8520), .a(n5658), .b(n7844), .c(net_253) );
ao22f01  g3033 ( .o(n8521), .a(n7847), .b(x4587), .c(n7846), .d(net_9815) );
na02f01  g3034 ( .o(n1464), .a(n8521), .b(n8520) );
no02f01  g3035 ( .o(n8523), .a(_net_9733), .b(_net_10157) );
in01f01  g3036 ( .o(n8524_1), .a(n8523) );
in01f01  g3037 ( .o(n8525), .a(_net_9733) );
no02f01  g3038 ( .o(n8526), .a(n8525), .b(n7797) );
ao12f01  g3039 ( .o(n8527), .a(n8526), .b(n8524_1), .c(n8134) );
in01f01  g3040 ( .o(n8528), .a(n8527) );
no02f01  g3041 ( .o(n8529_1), .a(n8135_1), .b(n8133) );
ao12f01  g3042 ( .o(n8530), .a(n8528), .b(n8529_1), .c(n8524_1) );
in01f01  g3043 ( .o(n8531), .a(n8530) );
in01f01  g3044 ( .o(n8532), .a(_net_9734) );
no02f01  g3045 ( .o(n8533), .a(n8532), .b(n7794) );
no02f01  g3046 ( .o(n8534_1), .a(_net_9734), .b(_net_10158) );
no02f01  g3047 ( .o(n8535), .a(n8534_1), .b(n8533) );
ao12f01  g3048 ( .o(n8536), .a(n6746), .b(n8535), .c(n8531) );
oa12f01  g3049 ( .o(n8537), .a(n8536), .b(n8535), .c(n8531) );
no02f01  g3050 ( .o(n8538_1), .a(n8145_1), .b(_net_10157) );
in01f01  g3051 ( .o(n8539), .a(n8538_1) );
no02f01  g3052 ( .o(n8540), .a(n8539), .b(_net_10158) );
in01f01  g3053 ( .o(n8541), .a(n8540) );
na02f01  g3054 ( .o(n8542), .a(n8539), .b(_net_10158) );
na02f01  g3055 ( .o(n8543_1), .a(n8542), .b(n8541) );
ao22f01  g3056 ( .o(n8544), .a(n8543_1), .b(n6750), .c(n6760), .d(_net_10158) );
na02f01  g3057 ( .o(n1469), .a(n8544), .b(n8537) );
na03f01  g3058 ( .o(n8546), .a(_net_9217), .b(n8089), .c(net_9216) );
in01f01  g3059 ( .o(n8547), .a(net_9210) );
na04f01  g3060 ( .o(n8548_1), .a(n8085), .b(n8547), .c(_net_9213), .d(n6672) );
no03f01  g3061 ( .o(n1478), .a(n8548_1), .b(n8546), .c(n8092) );
ao12f01  g3062 ( .o(n8550), .a(n5658), .b(n7844), .c(net_252) );
ao22f01  g3063 ( .o(n8551), .a(n7847), .b(x4694), .c(n7846), .d(net_9814) );
na02f01  g3064 ( .o(n1483), .a(n8551), .b(n8550) );
ao22f01  g3065 ( .o(n8553_1), .a(n5842), .b(net_9662), .c(n5841), .d(net_100) );
na02f01  g3066 ( .o(n8554), .a(n5847), .b(net_9959) );
ao22f01  g3067 ( .o(n8555), .a(n5850), .b(net_9761), .c(n5849_1), .d(net_9860) );
na03f01  g3068 ( .o(n1492), .a(n8555), .b(n8554), .c(n8553_1) );
in01f01  g3069 ( .o(n8557), .a(_net_9957) );
in01f01  g3070 ( .o(n8558_1), .a(_net_9958) );
na02f01  g3071 ( .o(n1497), .a(n8558_1), .b(n8557) );
in01f01  g3072 ( .o(n8560), .a(net_9848) );
oa22f01  g3073 ( .o(n1502), .a(n7480_1), .b(n8560), .c(n7478), .d(n5597_1) );
na02f01  g3074 ( .o(n8562_1), .a(n7782_1), .b(_net_10114) );
na02f01  g3075 ( .o(n1507), .a(n8562_1), .b(n7784) );
no02f01  g3076 ( .o(n8564), .a(n8161), .b(n8158) );
in01f01  g3077 ( .o(n8565), .a(n8564) );
ao12f01  g3078 ( .o(n8566), .a(n8184), .b(n8565), .c(n8174) );
oa12f01  g3079 ( .o(n8567_1), .a(n8566), .b(n8565), .c(n8174) );
na02f01  g3080 ( .o(n8568), .a(n8190_1), .b(_net_10366) );
na02f01  g3081 ( .o(n8569), .a(n8568), .b(n8192) );
ao22f01  g3082 ( .o(n8570), .a(n8569), .b(n8200_1), .c(n8202), .d(_net_10366) );
na02f01  g3083 ( .o(n1512), .a(n8570), .b(n8567_1) );
ao12f01  g3084 ( .o(n8572_1), .a(n5658), .b(n5678), .c(_net_259) );
ao22f01  g3085 ( .o(n8573), .a(n5681_1), .b(x4117), .c(n5680), .d(net_9722) );
na02f01  g3086 ( .o(n1526), .a(n8573), .b(n8572_1) );
in01f01  g3087 ( .o(n8575), .a(net_10193) );
in01f01  g3088 ( .o(n8576), .a(net_10188) );
na02f01  g3089 ( .o(n8577_1), .a(n8576), .b(x6599) );
in01f01  g3090 ( .o(n8578), .a(net_9568) );
in01f01  g3091 ( .o(n8579), .a(_net_9645) );
no04f01  g3092 ( .o(n8580), .a(n6009_1), .b(_net_9566), .c(n8579), .d(n8578) );
na02f01  g3093 ( .o(n8581), .a(n8580), .b(net_10175) );
ao12f01  g3094 ( .o(n1531), .a(n8577_1), .b(n8581), .c(n8575) );
in01f01  g3095 ( .o(n8583), .a(net_9825) );
na03f01  g3096 ( .o(n8584), .a(n8583), .b(n6801_1), .c(n6178) );
in01f01  g3097 ( .o(n8585), .a(net_9826) );
na04f01  g3098 ( .o(n8586), .a(n6773_1), .b(n6183), .c(n8585), .d(n6778_1) );
na04f01  g3099 ( .o(n8587_1), .a(n6904), .b(n6799), .c(n6785), .d(n6776) );
no03f01  g3100 ( .o(n8588), .a(n8587_1), .b(n8586), .c(n8584) );
ao12f01  g3101 ( .o(n1540), .a(n8588), .b(n6825), .c(n6769) );
ao12f01  g3102 ( .o(n8590), .a(n5658), .b(n5774), .c(x4285) );
oa12f01  g3103 ( .o(n1549), .a(n8590), .b(n5770), .c(n7048_1) );
in01f01  g3104 ( .o(n8592_1), .a(net_9849) );
oa22f01  g3105 ( .o(n1554), .a(n7480_1), .b(n8592_1), .c(n7478), .d(n5567_1) );
ao22f01  g3106 ( .o(n8594), .a(n8047), .b(net_10067), .c(n6564), .d(net_10089) );
oa12f01  g3107 ( .o(n8595), .a(n8594), .b(n6563), .c(n7753_1) );
ao22f01  g3108 ( .o(n8596), .a(n6592), .b(net_10176), .c(n6580), .d(net_9817) );
ao22f01  g3109 ( .o(n8597_1), .a(n6577), .b(net_9686), .c(n6572), .d(net_10386) );
na02f01  g3110 ( .o(n8598), .a(n8597_1), .b(n8596) );
no02f01  g3111 ( .o(n8599), .a(n8598), .b(n8595) );
ao22f01  g3112 ( .o(n8600), .a(n6606), .b(net_9947), .c(n6597), .d(net_9749) );
ao22f01  g3113 ( .o(n8601), .a(n6585), .b(net_9718), .c(n6584_1), .d(net_9785) );
na02f01  g3114 ( .o(n8602_1), .a(n6555), .b(net_9983) );
na02f01  g3115 ( .o(n8603), .a(n6602), .b(net_10015) );
na02f01  g3116 ( .o(n8604), .a(n8603), .b(n8602_1) );
in01f01  g3117 ( .o(n8605), .a(net_10046) );
na02f01  g3118 ( .o(n8606), .a(n6573), .b(net_9884) );
oa12f01  g3119 ( .o(n8607_1), .a(n8606), .b(n6591), .c(n8605) );
in01f01  g3120 ( .o(n8608), .a(net_10491) );
oa22f01  g3121 ( .o(n8609), .a(n8299), .b(n8608), .c(n6600), .d(n8560) );
in01f01  g3122 ( .o(n8610), .a(net_10281) );
na02f01  g3123 ( .o(n8611), .a(n6582), .b(net_9916) );
oa12f01  g3124 ( .o(n8612_1), .a(n8611), .b(n8302), .c(n8610) );
no04f01  g3125 ( .o(n8613), .a(n8612_1), .b(n8609), .c(n8607_1), .d(n8604) );
na04f01  g3126 ( .o(n1559), .a(n8613), .b(n8601), .c(n8600), .d(n8599) );
oa22f01  g3127 ( .o(n1564), .a(n7480_1), .b(n8585), .c(n7478), .d(n5513_1) );
na02f01  g3128 ( .o(n8616_1), .a(n6056), .b(net_260) );
na02f01  g3129 ( .o(n8617), .a(n6055), .b(net_9988) );
ao22f01  g3130 ( .o(n8618), .a(n6062_1), .b(x4041), .c(n6060), .d(_net_10439) );
na04f01  g3131 ( .o(n1569), .a(n8618), .b(n8617), .c(n8616_1), .d(n6058) );
in01f01  g3132 ( .o(n8620), .a(net_10045) );
in01f01  g3133 ( .o(n8621_1), .a(net_10036) );
no02f01  g3134 ( .o(n8622), .a(n6973), .b(n8621_1) );
na03f01  g3135 ( .o(n8623), .a(n5904), .b(x4520), .c(x6599) );
no02f01  g3136 ( .o(n8624), .a(n8622), .b(n5904) );
na02f01  g3137 ( .o(n8625), .a(n8624), .b(x6599) );
oa12f01  g3138 ( .o(n1574), .a(n8623), .b(n8625), .c(n8620) );
ao12f01  g3139 ( .o(n8627), .a(n5658), .b(n5678), .c(net_245) );
ao22f01  g3140 ( .o(n8628), .a(n5681_1), .b(x5225), .c(n5680), .d(net_9708) );
na02f01  g3141 ( .o(n1587), .a(n8628), .b(n8627) );
in01f01  g3142 ( .o(n8630), .a(_net_10113) );
ao12f01  g3143 ( .o(n8631_1), .a(n5658), .b(n6160_1), .c(x4937) );
oa12f01  g3144 ( .o(n1592), .a(n8631_1), .b(n6159), .c(n8630) );
ao12f01  g3145 ( .o(n8633), .a(n5658), .b(n5774), .c(x4694) );
oa12f01  g3146 ( .o(n1597), .a(n8633), .b(n5770), .c(n7018) );
in01f01  g3147 ( .o(n8635), .a(net_10047) );
oa22f01  g3148 ( .o(n1609), .a(n5907), .b(n8635), .c(n5905), .d(n5567_1) );
in01f01  g3149 ( .o(n8637), .a(n7923) );
no02f01  g3150 ( .o(n8638), .a(n8637), .b(n7883) );
in01f01  g3151 ( .o(n8639), .a(_net_9319) );
no02f01  g3152 ( .o(n8640), .a(n8639), .b(_net_9320) );
no02f01  g3153 ( .o(n8641_1), .a(_net_9319), .b(n8332) );
no02f01  g3154 ( .o(n8642), .a(n8641_1), .b(n8640) );
in01f01  g3155 ( .o(n8643), .a(net_9158) );
no02f01  g3156 ( .o(n8644), .a(n8643), .b(net_9159) );
in01f01  g3157 ( .o(n8645), .a(net_9159) );
no02f01  g3158 ( .o(n8646_1), .a(net_9158), .b(n8645) );
no02f01  g3159 ( .o(n8647), .a(n8646_1), .b(n8644) );
na02f01  g3160 ( .o(n8648), .a(n8647), .b(n8642) );
in01f01  g3161 ( .o(n8649), .a(n8642) );
in01f01  g3162 ( .o(n8650_1), .a(n8647) );
na02f01  g3163 ( .o(n8651), .a(n8650_1), .b(n8649) );
na03f01  g3164 ( .o(n8652), .a(n8651), .b(n8648), .c(n8638) );
ao12f01  g3165 ( .o(n8653), .a(n7883), .b(n8637), .c(_net_9313) );
na02f01  g3166 ( .o(n1614), .a(n8653), .b(n8652) );
in01f01  g3167 ( .o(n8655_1), .a(_net_10217) );
ao12f01  g3168 ( .o(n8656), .a(n5658), .b(n6887), .c(x5003) );
oa12f01  g3169 ( .o(n1631), .a(n8656), .b(n6885_1), .c(n8655_1) );
in01f01  g3170 ( .o(n8658), .a(_net_9322) );
ao12f01  g3171 ( .o(n8659_1), .a(n7883), .b(n7923), .c(_net_9314) );
oa12f01  g3172 ( .o(n1636), .a(n8659_1), .b(n7925_1), .c(n8658) );
in01f01  g3173 ( .o(n8661), .a(_net_9736) );
oa22f01  g3174 ( .o(n1641), .a(n7367), .b(n8661), .c(n7365_1), .d(n5585_1) );
na02f01  g3175 ( .o(n8663), .a(n6056), .b(net_253) );
na02f01  g3176 ( .o(n8664_1), .a(n6055), .b(net_9981) );
ao22f01  g3177 ( .o(n8665), .a(n6062_1), .b(x4587), .c(n6060), .d(_net_10432) );
na04f01  g3178 ( .o(n1646), .a(n8665), .b(n8664_1), .c(n8663), .d(n6058) );
in01f01  g3179 ( .o(n8667), .a(net_10077) );
oa22f01  g3180 ( .o(n1651), .a(n6989_1), .b(n5537_1), .c(n6988), .d(n8667) );
na02f01  g3181 ( .o(n8669), .a(n7353), .b(x5498) );
na02f01  g3182 ( .o(n8670), .a(n7352), .b(net_9672) );
ao22f01  g3183 ( .o(n8671), .a(n7358), .b(net_241), .c(n7357), .d(_net_10105) );
na04f01  g3184 ( .o(n1656), .a(n8671), .b(n8670), .c(n8669), .d(n7355_1) );
in01f01  g3185 ( .o(n8673_1), .a(n6621) );
na02f01  g3186 ( .o(n8674), .a(n8673_1), .b(n6619_1) );
oa12f01  g3187 ( .o(n8675), .a(n8674), .b(n6631), .c(n6620) );
no02f01  g3188 ( .o(n8676), .a(n6631), .b(n6620) );
in01f01  g3189 ( .o(n8677), .a(n8674) );
na02f01  g3190 ( .o(n8678_1), .a(n8677), .b(n8676) );
na02f01  g3191 ( .o(n1666), .a(n8678_1), .b(n8675) );
oa12f01  g3192 ( .o(n8680), .a(n7111), .b(n7306), .c(n7275_1) );
na03f01  g3193 ( .o(n8681), .a(n7318), .b(n7317_1), .c(n7108_1) );
na03f01  g3194 ( .o(n8682), .a(n8681), .b(n8680), .c(n6148) );
ao12f01  g3195 ( .o(n8683_1), .a(n6131_1), .b(n6147), .c(net_9367) );
na02f01  g3196 ( .o(n1671), .a(n8683_1), .b(n8682) );
in01f01  g3197 ( .o(n8685), .a(net_9954) );
in01f01  g3198 ( .o(n8686), .a(_net_232) );
in01f01  g3199 ( .o(n8687), .a(net_10539) );
oa12f01  g3200 ( .o(n8688_1), .a(x6599), .b(n6872), .c(n8687) );
no02f01  g3201 ( .o(n8689), .a(n8687), .b(n5658) );
na02f01  g3202 ( .o(n8690), .a(n8689), .b(net_10385) );
oa22f01  g3203 ( .o(n1676), .a(n8690), .b(n8686), .c(n8688_1), .d(n8685) );
ao22f01  g3204 ( .o(n8692), .a(n8118), .b(x3194), .c(n8117), .d(_net_9390) );
oa12f01  g3205 ( .o(n1681), .a(n8692), .b(n8116_1), .c(n5737) );
in01f01  g3206 ( .o(n8694), .a(n7896) );
no02f01  g3207 ( .o(n8695), .a(n7921_1), .b(n8694) );
na02f01  g3208 ( .o(n8696), .a(n8695), .b(net_9153) );
oa12f01  g3209 ( .o(n1686), .a(n8696), .b(n8695), .c(n6355) );
ao22f01  g3210 ( .o(n8698), .a(n5842), .b(net_9669), .c(n5841), .d(net_107) );
na02f01  g3211 ( .o(n8699), .a(n5847), .b(net_9966) );
ao22f01  g3212 ( .o(n8700), .a(n5850), .b(net_9768), .c(n5849_1), .d(net_9867) );
na03f01  g3213 ( .o(n1691), .a(n8700), .b(n8699), .c(n8698) );
na02f01  g3214 ( .o(n8702_1), .a(net_9651), .b(net_9650) );
in01f01  g3215 ( .o(n8703), .a(n8702_1) );
na02f01  g3216 ( .o(n8704), .a(n8703), .b(net_9652) );
no03f01  g3217 ( .o(n8705), .a(n8704), .b(n8420), .c(n8422) );
no02f01  g3218 ( .o(n8706), .a(n8704), .b(n8420) );
no02f01  g3219 ( .o(n8707_1), .a(n8706), .b(net_9654) );
no03f01  g3220 ( .o(n1696), .a(n8707_1), .b(n8705), .c(net_9151) );
in01f01  g3221 ( .o(n8709), .a(_net_10307) );
ao12f01  g3222 ( .o(n8710), .a(n5658), .b(n5774), .c(x5961) );
oa12f01  g3223 ( .o(n1701), .a(n8710), .b(n5770), .c(n8709) );
ao12f01  g3224 ( .o(n8712_1), .a(n5658), .b(n7737), .c(net_9350) );
oa12f01  g3225 ( .o(n1706), .a(n8712_1), .b(n7736), .c(n8645) );
in01f01  g3226 ( .o(n8714), .a(n7895) );
na02f01  g3227 ( .o(n8715), .a(net_225), .b(n6355) );
na04f01  g3228 ( .o(n8716), .a(n8715), .b(n8714), .c(net_9310), .d(_net_280) );
no02f01  g3229 ( .o(n8717_1), .a(net_9306), .b(net_229) );
in01f01  g3230 ( .o(n8718), .a(net_229) );
no02f01  g3231 ( .o(n8719), .a(n6407), .b(n8718) );
no02f01  g3232 ( .o(n8720), .a(net_227), .b(net_9304) );
no02f01  g3233 ( .o(n8721), .a(n8044), .b(n6367) );
oa22f01  g3234 ( .o(n8722_1), .a(n8721), .b(n8720), .c(n8719), .d(n8717_1) );
no02f01  g3235 ( .o(n8723), .a(n8722_1), .b(n8716) );
na02f01  g3236 ( .o(n8724), .a(n8021), .b(n6514) );
in01f01  g3237 ( .o(n8725), .a(net_224) );
oa22f01  g3238 ( .o(n8726), .a(net_225), .b(n6355), .c(n8725), .d(_net_9301) );
ao12f01  g3239 ( .o(n8727_1), .a(n8726), .b(n8725), .c(_net_9301) );
no02f01  g3240 ( .o(n8728), .a(net_9305), .b(net_228) );
no02f01  g3241 ( .o(n8729), .a(n6387), .b(n8416) );
oa22f01  g3242 ( .o(n8730), .a(n8729), .b(n8728), .c(n7901), .d(n7892) );
oa22f01  g3243 ( .o(n8731), .a(n7917), .b(n7901), .c(n7904), .d(n7892) );
no02f01  g3244 ( .o(n8732_1), .a(net_226), .b(net_9303) );
in01f01  g3245 ( .o(n8733), .a(net_226) );
no02f01  g3246 ( .o(n8734), .a(n8733), .b(n6362) );
no02f01  g3247 ( .o(n8735), .a(net_9307), .b(net_230) );
in01f01  g3248 ( .o(n8736), .a(net_230) );
no02f01  g3249 ( .o(n8737_1), .a(n6373_1), .b(n8736) );
oa22f01  g3250 ( .o(n8738), .a(n8737_1), .b(n8735), .c(n8734), .d(n8732_1) );
oa22f01  g3251 ( .o(n8739), .a(n7917), .b(n7904), .c(n7892), .d(n6459) );
no04f01  g3252 ( .o(n8740), .a(n8739), .b(n8738), .c(n8731), .d(n8730) );
na04f01  g3253 ( .o(n8741), .a(n8740), .b(n8727_1), .c(n8724), .d(n8723) );
no02f01  g3254 ( .o(n2827), .a(n8741), .b(n5633) );
in01f01  g3255 ( .o(n8743), .a(n2827) );
in01f01  g3256 ( .o(n8744), .a(_net_9637) );
in01f01  g3257 ( .o(n8745), .a(n7964) );
no02f01  g3258 ( .o(n8746), .a(n3455), .b(n2439) );
ao12f01  g3259 ( .o(n8747_1), .a(_net_187), .b(n8746), .c(n5918) );
in01f01  g3260 ( .o(n8748), .a(n8747_1) );
na04f01  g3261 ( .o(n8749), .a(n8748), .b(n7974), .c(n7968), .d(n8745) );
no02f01  g3262 ( .o(n8750), .a(n7972_1), .b(n8744) );
in01f01  g3263 ( .o(n8751), .a(n8750) );
no04f01  g3264 ( .o(n8752_1), .a(n8751), .b(n8749), .c(n7966), .d(n8744) );
in01f01  g3265 ( .o(n8753), .a(_net_9641) );
no02f01  g3266 ( .o(n8754), .a(n7732), .b(_net_9160) );
no02f01  g3267 ( .o(n8752), .a(n8754), .b(n7884) );
in01f01  g3268 ( .o(n8756), .a(n8752) );
in01f01  g3269 ( .o(n8757_1), .a(_net_9317) );
in01f01  g3270 ( .o(n8758), .a(_net_9318) );
in01f01  g3271 ( .o(n8759), .a(_net_9323) );
na04f01  g3272 ( .o(n8760), .a(n8759), .b(_net_9314), .c(n8758), .d(n8757_1) );
na04f01  g3273 ( .o(n8761), .a(n8658), .b(_net_9313), .c(n8332), .d(n7882) );
in01f01  g3274 ( .o(n8762_1), .a(_net_9324) );
in01f01  g3275 ( .o(n8763), .a(_net_9321) );
no02f01  g3276 ( .o(n8764), .a(_net_9315), .b(_net_9316) );
na03f01  g3277 ( .o(n8765), .a(n8764), .b(n8763), .c(n8762_1) );
na04f01  g3278 ( .o(n8766), .a(_net_9326), .b(_net_9311), .c(n8333), .d(n8639) );
no04f01  g3279 ( .o(n8767_1), .a(n8766), .b(n8765), .c(n8761), .d(n8760) );
no02f01  g3280 ( .o(n8768), .a(n8767_1), .b(n8756) );
no03f01  g3281 ( .o(n8769), .a(n8768), .b(_net_9250), .c(_net_9649) );
na02f01  g3282 ( .o(n8770), .a(n8756), .b(_net_9637) );
ao12f01  g3283 ( .o(n8771), .a(n8753), .b(n8770), .c(n8769) );
in01f01  g3284 ( .o(n8772_1), .a(_net_9640) );
no02f01  g3285 ( .o(n8773), .a(n8714), .b(n6354) );
in01f01  g3286 ( .o(n8774), .a(n8773) );
ao12f01  g3287 ( .o(n8775), .a(net_9612), .b(n8774), .c(_net_9637) );
no02f01  g3288 ( .o(n8776), .a(net_9648), .b(net_9647) );
in01f01  g3289 ( .o(n8777_1), .a(n8776) );
no03f01  g3290 ( .o(n8778), .a(n8777_1), .b(_net_9611), .c(_net_9250) );
in01f01  g3291 ( .o(n8779), .a(n8778) );
na02f01  g3292 ( .o(n8780), .a(n8779), .b(_net_9643) );
in01f01  g3293 ( .o(n8781), .a(net_9279) );
na03f01  g3294 ( .o(n8782_1), .a(n8781), .b(_net_9639), .c(_net_9637) );
in01f01  g3295 ( .o(n8783), .a(_net_9646) );
in01f01  g3296 ( .o(n8784), .a(_net_9638) );
na03f01  g3297 ( .o(n8785), .a(n8784), .b(n8783), .c(x6599) );
ao12f01  g3298 ( .o(n8786), .a(n8785), .b(_net_9250), .c(_net_9642) );
na03f01  g3299 ( .o(n8787_1), .a(n8786), .b(n8782_1), .c(n8780) );
ao12f01  g3300 ( .o(n8788), .a(n8787_1), .b(n7972_1), .c(_net_9637) );
oa12f01  g3301 ( .o(n8789), .a(n8788), .b(n8775), .c(n8772_1) );
no03f01  g3302 ( .o(n8790), .a(n8789), .b(n8771), .c(n8752_1) );
na02f01  g3303 ( .o(n1711), .a(n8790), .b(n8743) );
oa22f01  g3304 ( .o(n1720), .a(n6989_1), .b(n5576), .c(n6988), .d(n6556_1) );
in01f01  g3305 ( .o(n8793), .a(_net_10440) );
ao12f01  g3306 ( .o(n8794), .a(n5658), .b(n6052_1), .c(x3949) );
oa12f01  g3307 ( .o(n1725), .a(n8794), .b(n6048), .c(n8793) );
ao12f01  g3308 ( .o(n8796_1), .a(n5658), .b(n6875_1), .c(_net_232) );
ao22f01  g3309 ( .o(n8797), .a(n6878), .b(x6028), .c(n6877), .d(net_9893) );
na02f01  g3310 ( .o(n1730), .a(n8797), .b(n8796_1) );
ao12f01  g3311 ( .o(n8799), .a(n5658), .b(n5678), .c(_net_232) );
ao22f01  g3312 ( .o(n8800_1), .a(n5681_1), .b(x6028), .c(n5680), .d(net_9695) );
na02f01  g3313 ( .o(n1739), .a(n8800_1), .b(n8799) );
ao12f01  g3314 ( .o(n8802), .a(n5658), .b(n7844), .c(net_239) );
ao22f01  g3315 ( .o(n8803), .a(n7847), .b(x5601), .c(n7846), .d(net_9801) );
na02f01  g3316 ( .o(n1744), .a(n8803), .b(n8802) );
in01f01  g3317 ( .o(n8805), .a(net_9510) );
ao22f01  g3318 ( .o(n8806), .a(n5743), .b(x1459), .c(n5742), .d(_net_9419) );
oa12f01  g3319 ( .o(n1749), .a(n8806), .b(n5741), .c(n8805) );
oa22f01  g3320 ( .o(n1754), .a(n7480_1), .b(n6183), .c(n7478), .d(n5621) );
no03f01  g3321 ( .o(n8809_1), .a(net_9513), .b(n5738), .c(n5658) );
in01f01  g3322 ( .o(n8810), .a(n8809_1) );
no02f01  g3323 ( .o(n8811), .a(n6025), .b(n7593) );
in01f01  g3324 ( .o(n8812), .a(n8811) );
no02f01  g3325 ( .o(n8813), .a(n8812), .b(n7571_1) );
in01f01  g3326 ( .o(n8814_1), .a(n8813) );
na02f01  g3327 ( .o(n8815), .a(n8812), .b(n7571_1) );
na02f01  g3328 ( .o(n8816), .a(n8815), .b(n8814_1) );
na03f01  g3329 ( .o(n8817), .a(n5853_1), .b(n5738), .c(x6599) );
oa22f01  g3330 ( .o(n1759), .a(n8817), .b(n7571_1), .c(n8816), .d(n8810) );
na02f01  g3331 ( .o(n8819_1), .a(n5759), .b(_net_10123) );
na02f01  g3332 ( .o(n1764), .a(n8819_1), .b(n5761) );
in01f01  g3333 ( .o(n8821), .a(net_10190) );
na02f01  g3334 ( .o(n8822), .a(n8768), .b(net_10175) );
ao12f01  g3335 ( .o(n1769), .a(n8577_1), .b(n8822), .c(n8821) );
in01f01  g3336 ( .o(n8824_1), .a(_net_9189) );
oa22f01  g3337 ( .o(n1779), .a(n8349_1), .b(n8028), .c(n8347), .d(n8824_1) );
in01f01  g3338 ( .o(n8826), .a(net_9951) );
in01f01  g3339 ( .o(n8827), .a(_net_233) );
in01f01  g3340 ( .o(n8828), .a(net_10540) );
oa12f01  g3341 ( .o(n8829_1), .a(x6599), .b(n8828), .c(n6872) );
no02f01  g3342 ( .o(n8830), .a(n8828), .b(n5658) );
na02f01  g3343 ( .o(n8831), .a(n8830), .b(net_10385) );
oa22f01  g3344 ( .o(n1787), .a(n8831), .b(n8827), .c(n8829_1), .d(n8826) );
na02f01  g3345 ( .o(n8833), .a(n6020), .b(n5987) );
oa12f01  g3346 ( .o(n1792), .a(n8833), .b(n6020), .c(n5983_1) );
in01f01  g3347 ( .o(n8835), .a(net_9253) );
no02f01  g3348 ( .o(n8836), .a(n5938), .b(n8835) );
na02f01  g3349 ( .o(n8837), .a(n5938), .b(n8835) );
in01f01  g3350 ( .o(n8838), .a(n8837) );
na02f01  g3351 ( .o(n8839_1), .a(n6024), .b(net_9252) );
na02f01  g3352 ( .o(n8840), .a(n5935_1), .b(_net_117) );
oa12f01  g3353 ( .o(n8841), .a(n8840), .b(n5935_1), .c(n5946) );
na02f01  g3354 ( .o(n8842), .a(n8841), .b(net_9251) );
no02f01  g3355 ( .o(n8843), .a(n6024), .b(net_9252) );
oa12f01  g3356 ( .o(n8844_1), .a(n8839_1), .b(n8843), .c(n8842) );
oa12f01  g3357 ( .o(n8845), .a(n8844_1), .b(n8838), .c(n8836) );
in01f01  g3358 ( .o(n8846), .a(n8836) );
in01f01  g3359 ( .o(n8847), .a(n8844_1) );
na03f01  g3360 ( .o(n8848), .a(n8847), .b(n8837), .c(n8846) );
na02f01  g3361 ( .o(n1797), .a(n8848), .b(n8845) );
ao12f01  g3362 ( .o(n8850), .a(n6131_1), .b(n6148), .c(net_9364) );
oa12f01  g3363 ( .o(n1802), .a(n8850), .b(n8101_1), .c(n7097) );
no02f01  g3364 ( .o(n8852), .a(n5961), .b(n7708) );
in01f01  g3365 ( .o(n8853_1), .a(_net_9258) );
in01f01  g3366 ( .o(n8854), .a(n8852) );
oa12f01  g3367 ( .o(n8855), .a(n8853_1), .b(n8854), .c(n5958) );
oa12f01  g3368 ( .o(n8856), .a(n8855), .b(n8852), .c(n6614_1) );
no02f01  g3369 ( .o(n8857_1), .a(n6614_1), .b(_net_9258) );
in01f01  g3370 ( .o(n8858), .a(n8857_1) );
no02f01  g3371 ( .o(n8859), .a(n6634_1), .b(net_9257) );
in01f01  g3372 ( .o(n8860), .a(net_9255) );
no02f01  g3373 ( .o(n8861), .a(n5965), .b(n8860) );
in01f01  g3374 ( .o(n8862_1), .a(net_9256) );
in01f01  g3375 ( .o(n8863), .a(n8861) );
oa12f01  g3376 ( .o(n8864), .a(n8862_1), .b(n8863), .c(n5968) );
oa12f01  g3377 ( .o(n8865), .a(n8864), .b(n8861), .c(n5976) );
no02f01  g3378 ( .o(n8866), .a(n8865), .b(n8859) );
no02f01  g3379 ( .o(n8867_1), .a(n7072), .b(net_9254) );
na02f01  g3380 ( .o(n8868), .a(n8844_1), .b(n8837) );
no02f01  g3381 ( .o(n8869), .a(n8868), .b(n8867_1) );
in01f01  g3382 ( .o(n8870), .a(net_9254) );
no02f01  g3383 ( .o(n8871), .a(n5941), .b(n8870) );
na02f01  g3384 ( .o(n8872_1), .a(n5941), .b(n8870) );
oa12f01  g3385 ( .o(n8873), .a(n8872_1), .b(n8871), .c(n8836) );
in01f01  g3386 ( .o(n8874), .a(n8873) );
no02f01  g3387 ( .o(n8875), .a(n8874), .b(n8869) );
no02f01  g3388 ( .o(n8876_1), .a(n5976), .b(net_9256) );
no02f01  g3389 ( .o(n8877), .a(n6617), .b(net_9255) );
no03f01  g3390 ( .o(n8878), .a(n8877), .b(n8876_1), .c(n8859) );
in01f01  g3391 ( .o(n8879), .a(n8878) );
no02f01  g3392 ( .o(n8880), .a(n8879), .b(n8875) );
oa12f01  g3393 ( .o(n8881), .a(n8858), .b(n8880), .c(n8866) );
no02f01  g3394 ( .o(n8882), .a(n6017), .b(net_9263) );
no02f01  g3395 ( .o(n8883), .a(n6011), .b(net_9262) );
no02f01  g3396 ( .o(n8884), .a(n5987), .b(net_9261) );
no02f01  g3397 ( .o(n8885), .a(n8884), .b(n8883) );
in01f01  g3398 ( .o(n8886), .a(n8885) );
no02f01  g3399 ( .o(n8887), .a(n5994), .b(net_9260) );
no02f01  g3400 ( .o(n8888), .a(n5998_1), .b(net_9259) );
no02f01  g3401 ( .o(n8889), .a(n8888), .b(n8887) );
in01f01  g3402 ( .o(n8890), .a(n8889) );
no02f01  g3403 ( .o(n8891), .a(n8890), .b(n8886) );
in01f01  g3404 ( .o(n8892), .a(n8891) );
no02f01  g3405 ( .o(n8893), .a(n8892), .b(n8882) );
in01f01  g3406 ( .o(n8894), .a(n8893) );
ao12f01  g3407 ( .o(n8895), .a(n8894), .b(n8881), .c(n8856) );
in01f01  g3408 ( .o(n8896), .a(net_9262) );
in01f01  g3409 ( .o(n8897), .a(n6011) );
in01f01  g3410 ( .o(n8898), .a(net_9261) );
no02f01  g3411 ( .o(n8899), .a(n5986), .b(n8898) );
no02f01  g3412 ( .o(n8900), .a(n8897), .b(n8896) );
no02f01  g3413 ( .o(n8901), .a(n8900), .b(n8899) );
ao12f01  g3414 ( .o(n8902), .a(n8901), .b(n8897), .c(n8896) );
in01f01  g3415 ( .o(n8903), .a(net_9259) );
no02f01  g3416 ( .o(n8904), .a(n5997), .b(n8903) );
in01f01  g3417 ( .o(n8905), .a(n8904) );
ao12f01  g3418 ( .o(n8906), .a(net_9260), .b(n8904), .c(n5994) );
ao12f01  g3419 ( .o(n8907), .a(n8906), .b(n8905), .c(n5993_1) );
ao12f01  g3420 ( .o(n8908), .a(n8902), .b(n8907), .c(n8885) );
no02f01  g3421 ( .o(n8909), .a(n8908), .b(n8882) );
in01f01  g3422 ( .o(n8910), .a(n8909) );
in01f01  g3423 ( .o(n8911), .a(net_9263) );
in01f01  g3424 ( .o(n8912), .a(n6017) );
no02f01  g3425 ( .o(n8913), .a(n8912), .b(n8911) );
in01f01  g3426 ( .o(n8914), .a(n8913) );
na02f01  g3427 ( .o(n8915), .a(n8914), .b(n8910) );
no02f01  g3428 ( .o(n8916), .a(n8915), .b(n8895) );
in01f01  g3429 ( .o(n8917), .a(net_9264) );
in01f01  g3430 ( .o(n8918), .a(n6014) );
no02f01  g3431 ( .o(n8919), .a(n8918), .b(n8917) );
no02f01  g3432 ( .o(n8920), .a(n6014), .b(net_9264) );
no02f01  g3433 ( .o(n8921), .a(n8920), .b(n8919) );
na02f01  g3434 ( .o(n8922), .a(n8921), .b(n8916) );
in01f01  g3435 ( .o(n8923), .a(n8921) );
oa12f01  g3436 ( .o(n8924), .a(n8923), .b(n8915), .c(n8895) );
na02f01  g3437 ( .o(n1807), .a(n8924), .b(n8922) );
ao12f01  g3438 ( .o(n8926), .a(n5658), .b(n6160_1), .c(x4781) );
oa12f01  g3439 ( .o(n1812), .a(n8926), .b(n6159), .c(n7780) );
no02f01  g3440 ( .o(n7695), .a(n6021), .b(n8912) );
in01f01  g3441 ( .o(n8929), .a(n7695) );
no02f01  g3442 ( .o(n1817), .a(n8929), .b(n5927) );
in01f01  g3443 ( .o(n8931), .a(_net_10335) );
no02f01  g3444 ( .o(n8932), .a(_net_10329), .b(_net_10328) );
in01f01  g3445 ( .o(n8933), .a(n8932) );
ao12f01  g3446 ( .o(n8934), .a(_net_10326), .b(_net_10325), .c(_net_10324) );
in01f01  g3447 ( .o(n8935), .a(n8934) );
no02f01  g3448 ( .o(n8936), .a(n8935), .b(_net_10327) );
in01f01  g3449 ( .o(n8937), .a(n8936) );
no02f01  g3450 ( .o(n8938), .a(n8937), .b(n8933) );
in01f01  g3451 ( .o(n8939), .a(n8938) );
no02f01  g3452 ( .o(n8940), .a(n8939), .b(_net_10330) );
in01f01  g3453 ( .o(n8941), .a(n8940) );
no02f01  g3454 ( .o(n8942), .a(n8941), .b(_net_10331) );
in01f01  g3455 ( .o(n8943), .a(n8942) );
no02f01  g3456 ( .o(n8944), .a(n8943), .b(_net_10332) );
in01f01  g3457 ( .o(n8945), .a(n8944) );
no02f01  g3458 ( .o(n8946), .a(n8945), .b(_net_10333) );
in01f01  g3459 ( .o(n8947), .a(n8946) );
no02f01  g3460 ( .o(n8948), .a(n8947), .b(_net_10334) );
na02f01  g3461 ( .o(n8949), .a(n8948), .b(n8931) );
in01f01  g3462 ( .o(n8950), .a(n8948) );
na02f01  g3463 ( .o(n8951), .a(n8950), .b(_net_10335) );
na02f01  g3464 ( .o(n1822), .a(n8951), .b(n8949) );
ao22f01  g3465 ( .o(n8953), .a(n5842), .b(net_9689), .c(n5841), .d(_net_127) );
na02f01  g3466 ( .o(n8954), .a(n5847), .b(net_9986) );
ao22f01  g3467 ( .o(n8955), .a(n5850), .b(net_9788), .c(n5849_1), .d(net_9887) );
na03f01  g3468 ( .o(n1835), .a(n8955), .b(n8954), .c(n8953) );
in01f01  g3469 ( .o(n8957), .a(_net_10221) );
no02f01  g3470 ( .o(n8958), .a(_net_10259), .b(n8957) );
no02f01  g3471 ( .o(n8959), .a(n6903), .b(_net_10221) );
in01f01  g3472 ( .o(n8960), .a(_net_10220) );
no02f01  g3473 ( .o(n8961), .a(n8960), .b(_net_10258) );
no02f01  g3474 ( .o(n8962), .a(n6172), .b(_net_10219) );
in01f01  g3475 ( .o(n8963), .a(n8962) );
no02f01  g3476 ( .o(n8964), .a(_net_10220), .b(n6171) );
in01f01  g3477 ( .o(n8965), .a(n8964) );
ao12f01  g3478 ( .o(n8966), .a(n8961), .b(n8965), .c(n8963) );
no02f01  g3479 ( .o(n8967), .a(n8966), .b(n8959) );
no02f01  g3480 ( .o(n8968), .a(_net_10222), .b(n6902) );
in01f01  g3481 ( .o(n8969), .a(_net_10222) );
no02f01  g3482 ( .o(n8970), .a(n8969), .b(_net_10260) );
no02f01  g3483 ( .o(n8971), .a(n8970), .b(n8968) );
in01f01  g3484 ( .o(n8972), .a(n8971) );
oa12f01  g3485 ( .o(n8973), .a(n8972), .b(n8967), .c(n8958) );
in01f01  g3486 ( .o(n8974), .a(n8958) );
in01f01  g3487 ( .o(n8975), .a(n8967) );
na03f01  g3488 ( .o(n8976), .a(n8971), .b(n8975), .c(n8974) );
na02f01  g3489 ( .o(n1844), .a(n8976), .b(n8973) );
in01f01  g3490 ( .o(n8978), .a(_net_10227) );
ao12f01  g3491 ( .o(n8979), .a(n5658), .b(n6887), .c(x4209) );
oa12f01  g3492 ( .o(n1849), .a(n8979), .b(n6885_1), .c(n8978) );
no02f01  g3493 ( .o(n8981), .a(n8762_1), .b(_net_9323) );
no02f01  g3494 ( .o(n8982), .a(_net_9324), .b(n8759) );
no02f01  g3495 ( .o(n8983), .a(n8982), .b(n8981) );
in01f01  g3496 ( .o(n8984), .a(net_9154) );
no02f01  g3497 ( .o(n8985), .a(net_9155), .b(n8984) );
no02f01  g3498 ( .o(n8986), .a(n7731), .b(net_9154) );
no02f01  g3499 ( .o(n8987), .a(n8986), .b(n8985) );
na02f01  g3500 ( .o(n8988), .a(n8987), .b(n8983) );
in01f01  g3501 ( .o(n8989), .a(n8983) );
in01f01  g3502 ( .o(n8990), .a(n8987) );
na02f01  g3503 ( .o(n8991), .a(n8990), .b(n8989) );
na03f01  g3504 ( .o(n8992), .a(n8991), .b(n8988), .c(n8638) );
ao12f01  g3505 ( .o(n8993), .a(n7883), .b(n8637), .c(_net_9317) );
na02f01  g3506 ( .o(n1854), .a(n8993), .b(n8992) );
in01f01  g3507 ( .o(n8995), .a(net_9738) );
oa22f01  g3508 ( .o(n1859), .a(n7367), .b(n8995), .c(n7365_1), .d(n5634) );
ao22f01  g3509 ( .o(n8997), .a(n5842), .b(net_9717), .c(n5841), .d(_net_157) );
na02f01  g3510 ( .o(n8998), .a(n5847), .b(net_10014) );
ao22f01  g3511 ( .o(n8999), .a(n5850), .b(net_9816), .c(n5849_1), .d(net_9915) );
na03f01  g3512 ( .o(n1868), .a(n8999), .b(n8998), .c(n8997) );
ao12f01  g3513 ( .o(n9001), .a(n5658), .b(n6532), .c(net_260) );
ao22f01  g3514 ( .o(n9002), .a(n6535), .b(x4041), .c(n6534), .d(net_10020) );
na02f01  g3515 ( .o(n1877), .a(n9002), .b(n9001) );
no03f01  g3516 ( .o(n9004), .a(_net_10477), .b(_net_10476), .c(_net_10475) );
na03f01  g3517 ( .o(n9005), .a(n9004), .b(n7433), .c(n7369) );
no04f01  g3518 ( .o(n9006), .a(_net_10472), .b(_net_10474), .c(_net_10471), .d(_net_10473) );
na02f01  g3519 ( .o(n9007), .a(n9006), .b(n7436_1) );
no02f01  g3520 ( .o(n9008), .a(n9007), .b(n9005) );
in01f01  g3521 ( .o(n9009), .a(_net_10049) );
no02f01  g3522 ( .o(n9010), .a(n9009), .b(_net_10048) );
in01f01  g3523 ( .o(n9011), .a(n9010) );
no03f01  g3524 ( .o(n9012), .a(n9011), .b(n9008), .c(n7429) );
in01f01  g3525 ( .o(n9013), .a(_net_10456) );
in01f01  g3526 ( .o(n9014), .a(_net_10455) );
ao22f01  g3527 ( .o(n9015), .a(n9014), .b(_net_10429), .c(n9013), .d(_net_10430) );
no02f01  g3528 ( .o(n9016), .a(n9015), .b(_net_10456) );
in01f01  g3529 ( .o(n9017), .a(_net_10458) );
in01f01  g3530 ( .o(n9018), .a(_net_10457) );
ao22f01  g3531 ( .o(n9019), .a(_net_10432), .b(n9017), .c(n9018), .d(_net_10431) );
oa12f01  g3532 ( .o(n9020), .a(n9019), .b(n9015), .c(n8227_1) );
ao12f01  g3533 ( .o(n9021), .a(n9018), .b(_net_10432), .c(n9017) );
ao22f01  g3534 ( .o(n9022), .a(n9021), .b(n7361), .c(n8219_1), .d(_net_10458) );
oa12f01  g3535 ( .o(n9023), .a(n9022), .b(n9020), .c(n9016) );
in01f01  g3536 ( .o(n9024), .a(_net_10460) );
in01f01  g3537 ( .o(n9025), .a(_net_10459) );
ao22f01  g3538 ( .o(n9026), .a(n9025), .b(_net_10433), .c(n9024), .d(_net_10434) );
in01f01  g3539 ( .o(n9027), .a(_net_10436) );
oa22f01  g3540 ( .o(n9028), .a(_net_10462), .b(n9027), .c(_net_10461), .d(n8240_1) );
in01f01  g3541 ( .o(n9029), .a(n9028) );
na03f01  g3542 ( .o(n9030), .a(n9029), .b(n9026), .c(n9023) );
na03f01  g3543 ( .o(n9031), .a(n9029), .b(_net_10460), .c(n8209) );
no02f01  g3544 ( .o(n9032), .a(n9025), .b(n9024) );
in01f01  g3545 ( .o(n9033), .a(n9032) );
oa22f01  g3546 ( .o(n9034), .a(n9033), .b(_net_10433), .c(n7664), .d(n9025) );
na02f01  g3547 ( .o(n9035), .a(n9034), .b(n9029) );
in01f01  g3548 ( .o(n9036), .a(_net_10461) );
in01f01  g3549 ( .o(n9037), .a(_net_10462) );
ao12f01  g3550 ( .o(n9038), .a(n9036), .b(n9037), .c(_net_10436) );
ao22f01  g3551 ( .o(n9039), .a(n9038), .b(n8240_1), .c(_net_10462), .d(n9027) );
na04f01  g3552 ( .o(n9040), .a(n9039), .b(n9035), .c(n9031), .d(n9030) );
in01f01  g3553 ( .o(n9041), .a(_net_10439) );
oa22f01  g3554 ( .o(n9042), .a(_net_10466), .b(n8793), .c(n9041), .d(_net_10465) );
in01f01  g3555 ( .o(n9043), .a(_net_10438) );
in01f01  g3556 ( .o(n9044), .a(_net_10437) );
oa22f01  g3557 ( .o(n9045), .a(n9044), .b(_net_10463), .c(n9043), .d(_net_10464) );
no02f01  g3558 ( .o(n9046), .a(n9045), .b(n9042) );
na02f01  g3559 ( .o(n9047), .a(n9046), .b(n9040) );
in01f01  g3560 ( .o(n9048), .a(_net_10464) );
no03f01  g3561 ( .o(n9049), .a(n9042), .b(_net_10438), .c(n9048) );
oa12f01  g3562 ( .o(n9050), .a(_net_10463), .b(n9043), .c(_net_10464) );
no03f01  g3563 ( .o(n9051), .a(n9050), .b(n9042), .c(_net_10437) );
oa12f01  g3564 ( .o(n9052), .a(_net_10465), .b(_net_10466), .c(n8793) );
no02f01  g3565 ( .o(n9053), .a(n9052), .b(_net_10439) );
in01f01  g3566 ( .o(n9054), .a(_net_10466) );
in01f01  g3567 ( .o(n9055), .a(_net_10048) );
no03f01  g3568 ( .o(n9056), .a(_net_10049), .b(n7429), .c(n9055) );
oa12f01  g3569 ( .o(n9057), .a(n9056), .b(n9054), .c(_net_10440) );
no04f01  g3570 ( .o(n9058), .a(n9057), .b(n9053), .c(n9051), .d(n9049) );
ao12f01  g3571 ( .o(n9059), .a(n9012), .b(n9058), .c(n9047) );
no04f01  g3572 ( .o(n1886), .a(n9059), .b(net_10513), .c(net_10514), .d(_net_10512) );
no02f01  g3573 ( .o(n9061), .a(_net_10223), .b(_net_10224) );
in01f01  g3574 ( .o(n9062), .a(n9061) );
ao12f01  g3575 ( .o(n9063), .a(_net_10221), .b(_net_10220), .c(_net_10219) );
in01f01  g3576 ( .o(n9064), .a(n9063) );
no02f01  g3577 ( .o(n9065), .a(n9064), .b(_net_10222) );
in01f01  g3578 ( .o(n9066), .a(n9065) );
no02f01  g3579 ( .o(n9067), .a(n9066), .b(n9062) );
in01f01  g3580 ( .o(n9068), .a(n9067) );
no02f01  g3581 ( .o(n9069), .a(n9068), .b(_net_10225) );
in01f01  g3582 ( .o(n9070), .a(n9069) );
no02f01  g3583 ( .o(n9071), .a(n9070), .b(_net_10226) );
in01f01  g3584 ( .o(n9072), .a(n9071) );
no02f01  g3585 ( .o(n9073), .a(n9072), .b(_net_10227) );
in01f01  g3586 ( .o(n9074), .a(n9073) );
na02f01  g3587 ( .o(n9075), .a(n9072), .b(_net_10227) );
na02f01  g3588 ( .o(n1891), .a(n9075), .b(n9074) );
in01f01  g3589 ( .o(n9077), .a(_net_10359) );
in01f01  g3590 ( .o(n9078), .a(_net_10358) );
no02f01  g3591 ( .o(n9079), .a(_net_9934), .b(n9078) );
no02f01  g3592 ( .o(n9080), .a(n5705_1), .b(_net_10358) );
in01f01  g3593 ( .o(n9081), .a(n9080) );
no02f01  g3594 ( .o(n9082), .a(n5719_1), .b(_net_10357) );
no02f01  g3595 ( .o(n9083), .a(_net_10356), .b(n5718) );
no02f01  g3596 ( .o(n9084), .a(n5722), .b(_net_10355) );
in01f01  g3597 ( .o(n9085), .a(n9084) );
no02f01  g3598 ( .o(n9086), .a(_net_10354), .b(n5721) );
in01f01  g3599 ( .o(n9087), .a(_net_10352) );
no02f01  g3600 ( .o(n9088), .a(_net_9928), .b(n9087) );
in01f01  g3601 ( .o(n9089), .a(_net_10353) );
no02f01  g3602 ( .o(n9090), .a(n9089), .b(_net_9929) );
no02f01  g3603 ( .o(n9091), .a(n9090), .b(n9088) );
in01f01  g3604 ( .o(n9092), .a(n9091) );
no02f01  g3605 ( .o(n9093), .a(n5711), .b(_net_10352) );
na02f01  g3606 ( .o(n9094), .a(n5706), .b(_net_10351) );
no02f01  g3607 ( .o(n9095), .a(n5707), .b(_net_10350) );
no02f01  g3608 ( .o(n9096), .a(n5706), .b(_net_10351) );
oa12f01  g3609 ( .o(n9097), .a(n9094), .b(n9096), .c(n9095) );
in01f01  g3610 ( .o(n9098), .a(n9097) );
no02f01  g3611 ( .o(n9099), .a(n9098), .b(n9093) );
oa22f01  g3612 ( .o(n9100), .a(n9099), .b(n9092), .c(_net_10353), .d(n5710_1) );
no02f01  g3613 ( .o(n9101), .a(n9100), .b(n9086) );
na02f01  g3614 ( .o(n9102), .a(n9101), .b(n9085) );
no02f01  g3615 ( .o(n9103), .a(n9102), .b(n9083) );
in01f01  g3616 ( .o(n9104), .a(_net_10355) );
no02f01  g3617 ( .o(n9105), .a(_net_9931), .b(n9104) );
in01f01  g3618 ( .o(n9106), .a(_net_10354) );
no02f01  g3619 ( .o(n9107), .a(n9106), .b(_net_9930) );
ao12f01  g3620 ( .o(n9108), .a(n9105), .b(n9107), .c(n9085) );
no02f01  g3621 ( .o(n9109), .a(n9108), .b(n9083) );
in01f01  g3622 ( .o(n9110), .a(_net_10356) );
no02f01  g3623 ( .o(n9111), .a(n9110), .b(_net_9932) );
in01f01  g3624 ( .o(n9112), .a(_net_10357) );
no02f01  g3625 ( .o(n9113), .a(_net_9933), .b(n9112) );
no02f01  g3626 ( .o(n9114), .a(n9113), .b(n9111) );
ao12f01  g3627 ( .o(n9115), .a(n9114), .b(n9082), .c(_net_9933) );
no02f01  g3628 ( .o(n9116), .a(n9115), .b(n9109) );
in01f01  g3629 ( .o(n9117), .a(n9116) );
no02f01  g3630 ( .o(n9118), .a(n9117), .b(n9103) );
na02f01  g3631 ( .o(n9119), .a(n9115), .b(_net_10357) );
oa12f01  g3632 ( .o(n9120), .a(n9119), .b(n9118), .c(n9082) );
ao12f01  g3633 ( .o(n9121), .a(n9079), .b(n9120), .c(n9081) );
na02f01  g3634 ( .o(n9122), .a(n9121), .b(n9077) );
in01f01  g3635 ( .o(n9123), .a(n9122) );
no02f01  g3636 ( .o(n9124), .a(n9121), .b(n9077) );
oa12f01  g3637 ( .o(n9125), .a(n8183), .b(n9124), .c(n9123) );
no02f01  g3638 ( .o(n9126), .a(n9106), .b(n9104) );
in01f01  g3639 ( .o(n9127), .a(n9126) );
in01f01  g3640 ( .o(n9128), .a(_net_10351) );
in01f01  g3641 ( .o(n9129), .a(_net_10350) );
no02f01  g3642 ( .o(n9130), .a(n9129), .b(n9128) );
in01f01  g3643 ( .o(n9131), .a(n9130) );
no02f01  g3644 ( .o(n9132), .a(n9131), .b(n9087) );
in01f01  g3645 ( .o(n9133), .a(n9132) );
no02f01  g3646 ( .o(n9134), .a(n9133), .b(n9089) );
in01f01  g3647 ( .o(n9135), .a(n9134) );
no02f01  g3648 ( .o(n9136), .a(n9135), .b(n9127) );
in01f01  g3649 ( .o(n9137), .a(n9136) );
no02f01  g3650 ( .o(n9138), .a(n9137), .b(n9110) );
in01f01  g3651 ( .o(n9139), .a(n9138) );
no02f01  g3652 ( .o(n9140), .a(n9139), .b(n9112) );
na02f01  g3653 ( .o(n9141), .a(n9140), .b(_net_10358) );
no02f01  g3654 ( .o(n9142), .a(n9141), .b(n9077) );
in01f01  g3655 ( .o(n9143), .a(n9142) );
in01f01  g3656 ( .o(n9144), .a(n8200_1) );
ao12f01  g3657 ( .o(n9145), .a(n9144), .b(n9141), .c(n9077) );
ao22f01  g3658 ( .o(n9146), .a(n9145), .b(n9143), .c(n8202), .d(_net_10359) );
na02f01  g3659 ( .o(n1896), .a(n9146), .b(n9125) );
na02f01  g3660 ( .o(n9148), .a(n6349), .b(n6280) );
oa22f01  g3661 ( .o(n1901), .a(n9148), .b(n6348), .c(n6349), .d(n8862_1) );
in01f01  g3662 ( .o(n9150), .a(n6628) );
in01f01  g3663 ( .o(n9151), .a(n6629_1) );
no02f01  g3664 ( .o(n9152), .a(n9151), .b(n9150) );
oa22f01  g3665 ( .o(n9153), .a(n9152), .b(n6627), .c(n6626), .d(n6620) );
no02f01  g3666 ( .o(n9154), .a(n6626), .b(n6620) );
na02f01  g3667 ( .o(n9155), .a(n9154), .b(n6630) );
na02f01  g3668 ( .o(n1906), .a(n9155), .b(n9153) );
oa12f01  g3669 ( .o(n9157), .a(n6349), .b(n6271), .c(n6270) );
oa22f01  g3670 ( .o(n1911), .a(n9157), .b(n6348), .c(n6349), .d(n8835) );
in01f01  g3671 ( .o(n9159), .a(net_9289) );
na02f01  g3672 ( .o(n9160), .a(n6136_1), .b(_net_9380) );
ao12f01  g3673 ( .o(n1916), .a(n5658), .b(n9160), .c(n9159) );
in01f01  g3674 ( .o(n9162), .a(net_10497) );
oa22f01  g3675 ( .o(n1921), .a(n7467), .b(n5576), .c(n7465_1), .d(n9162) );
ao22f01  g3676 ( .o(n9164), .a(n5842), .b(_net_9751), .c(n5841), .d(_net_187) );
na02f01  g3677 ( .o(n9165), .a(n5847), .b(_net_10048) );
ao22f01  g3678 ( .o(n9166), .a(n5850), .b(_net_9850), .c(n5849_1), .d(_net_9949) );
na03f01  g3679 ( .o(n1926), .a(n9166), .b(n9165), .c(n9164) );
in01f01  g3680 ( .o(n9168), .a(net_9156) );
ao12f01  g3681 ( .o(n9169), .a(n5658), .b(n7737), .c(net_9347) );
oa12f01  g3682 ( .o(n1931), .a(n9169), .b(n7736), .c(n9168) );
in01f01  g3683 ( .o(n9171), .a(_net_10267) );
in01f01  g3684 ( .o(n9172), .a(_net_10228) );
no02f01  g3685 ( .o(n9173), .a(_net_10266), .b(n9172) );
in01f01  g3686 ( .o(n9174), .a(n9173) );
in01f01  g3687 ( .o(n9175), .a(_net_10266) );
no02f01  g3688 ( .o(n9176), .a(n9175), .b(_net_10228) );
no02f01  g3689 ( .o(n9177), .a(_net_10265), .b(n8978) );
in01f01  g3690 ( .o(n9178), .a(n9177) );
oa12f01  g3691 ( .o(n9179), .a(n9174), .b(n9178), .c(n9176) );
in01f01  g3692 ( .o(n9180), .a(_net_10229) );
in01f01  g3693 ( .o(n9181), .a(n9179) );
oa12f01  g3694 ( .o(n9182), .a(n9180), .b(n9181), .c(_net_10267) );
oa12f01  g3695 ( .o(n9183), .a(n9182), .b(n9179), .c(n9171) );
in01f01  g3696 ( .o(n9184), .a(n9183) );
in01f01  g3697 ( .o(n9185), .a(_net_10265) );
no02f01  g3698 ( .o(n9186), .a(n9185), .b(_net_10227) );
no02f01  g3699 ( .o(n9187), .a(_net_10226), .b(n6928) );
no02f01  g3700 ( .o(n9188), .a(_net_10223), .b(n6918) );
no02f01  g3701 ( .o(n9189), .a(n8970), .b(n8958) );
ao22f01  g3702 ( .o(n9190), .a(n9189), .b(n8975), .c(n8969), .d(_net_10260) );
in01f01  g3703 ( .o(n9191), .a(n9190) );
no02f01  g3704 ( .o(n9192), .a(n9191), .b(n9188) );
no02f01  g3705 ( .o(n9193), .a(n6923), .b(_net_10225) );
in01f01  g3706 ( .o(n9194), .a(n9193) );
no02f01  g3707 ( .o(n9195), .a(n6916), .b(_net_10224) );
in01f01  g3708 ( .o(n9196), .a(n9195) );
na03f01  g3709 ( .o(n9197), .a(n9196), .b(n9194), .c(n9192) );
in01f01  g3710 ( .o(n9198), .a(_net_10224) );
no02f01  g3711 ( .o(n9199), .a(_net_10262), .b(n9198) );
in01f01  g3712 ( .o(n9200), .a(_net_10223) );
no02f01  g3713 ( .o(n9201), .a(n9200), .b(_net_10261) );
ao12f01  g3714 ( .o(n9202), .a(n9199), .b(n9201), .c(n9196) );
no02f01  g3715 ( .o(n9203), .a(n9202), .b(n9193) );
in01f01  g3716 ( .o(n9204), .a(_net_10226) );
in01f01  g3717 ( .o(n9205), .a(_net_10225) );
no02f01  g3718 ( .o(n9206), .a(_net_10263), .b(n9205) );
no02f01  g3719 ( .o(n9207), .a(n9204), .b(_net_10264) );
no02f01  g3720 ( .o(n9208), .a(n9207), .b(n9206) );
ao12f01  g3721 ( .o(n9209), .a(n9208), .b(n9187), .c(n9204) );
no02f01  g3722 ( .o(n9210), .a(n9209), .b(n9203) );
ao12f01  g3723 ( .o(n9211), .a(n9187), .b(n9210), .c(n9197) );
na02f01  g3724 ( .o(n9212), .a(n9209), .b(n6928) );
in01f01  g3725 ( .o(n9213), .a(n9212) );
no02f01  g3726 ( .o(n9214), .a(n9213), .b(n9211) );
no02f01  g3727 ( .o(n9215), .a(n9214), .b(n9186) );
no02f01  g3728 ( .o(n9216), .a(n9171), .b(_net_10229) );
no02f01  g3729 ( .o(n9217), .a(n9216), .b(n9176) );
ao12f01  g3730 ( .o(n9218), .a(n9184), .b(n9217), .c(n9215) );
in01f01  g3731 ( .o(n9219), .a(n9218) );
in01f01  g3732 ( .o(n9220), .a(_net_10230) );
in01f01  g3733 ( .o(n9221), .a(_net_10268) );
no02f01  g3734 ( .o(n9222), .a(n9221), .b(n9220) );
no02f01  g3735 ( .o(n9223), .a(_net_10268), .b(_net_10230) );
no02f01  g3736 ( .o(n9224), .a(n9223), .b(n9222) );
na02f01  g3737 ( .o(n9225), .a(n9224), .b(n9219) );
in01f01  g3738 ( .o(n9226), .a(n9224) );
na02f01  g3739 ( .o(n9227), .a(n9226), .b(n9218) );
na02f01  g3740 ( .o(n1936), .a(n9227), .b(n9225) );
in01f01  g3741 ( .o(n9229), .a(_net_10231) );
ao12f01  g3742 ( .o(n9230), .a(n5658), .b(n6887), .c(x3889) );
oa12f01  g3743 ( .o(n1941), .a(n9230), .b(n6885_1), .c(n9229) );
in01f01  g3744 ( .o(n9232), .a(net_10493) );
oa22f01  g3745 ( .o(n1946), .a(n7467), .b(n5609), .c(n7465_1), .d(n9232) );
in01f01  g3746 ( .o(n9234), .a(_net_10420) );
ao12f01  g3747 ( .o(n9235), .a(n5658), .b(n6052_1), .c(x5498) );
oa12f01  g3748 ( .o(n1951), .a(n9235), .b(n6048), .c(n9234) );
in01f01  g3749 ( .o(n9237), .a(net_211) );
in01f01  g3750 ( .o(n9238), .a(net_10083) );
oa22f01  g3751 ( .o(n9239), .a(n6565), .b(n9238), .c(n6563), .d(n9237) );
ao12f01  g3752 ( .o(n9240), .a(n9239), .b(n6555), .c(net_9977) );
ao22f01  g3753 ( .o(n9241), .a(n6573), .b(net_9878), .c(n6572), .d(net_10394) );
ao22f01  g3754 ( .o(n9242), .a(n6580), .b(net_9811), .c(n6577), .d(net_9680) );
na02f01  g3755 ( .o(n9243), .a(n6584_1), .b(net_9779) );
ao22f01  g3756 ( .o(n9244), .a(n6599_1), .b(_net_9842), .c(n6582), .d(net_9910) );
na02f01  g3757 ( .o(n9245), .a(n9244), .b(n9243) );
ao22f01  g3758 ( .o(n9246), .a(n6592), .b(net_10184), .c(n6590), .d(_net_10040) );
ao22f01  g3759 ( .o(n9247), .a(n6597), .b(_net_9743), .c(n6585), .d(net_9712) );
ao22f01  g3760 ( .o(n9248), .a(n6603), .b(net_10499), .c(n6602), .d(net_10009) );
ao22f01  g3761 ( .o(n9249), .a(n6606), .b(_net_9941), .c(n6605), .d(net_10289) );
na04f01  g3762 ( .o(n9250), .a(n9249), .b(n9248), .c(n9247), .d(n9246) );
no02f01  g3763 ( .o(n9251), .a(n9250), .b(n9245) );
na04f01  g3764 ( .o(n1956), .a(n9251), .b(n9242), .c(n9241), .d(n9240) );
in01f01  g3765 ( .o(n9253), .a(net_10178) );
oa22f01  g3766 ( .o(n1960), .a(n7956), .b(n5609), .c(n7955), .d(n9253) );
no04f01  g3767 ( .o(n9255), .a(n8179), .b(n8174), .c(n8161), .d(n8155_1) );
in01f01  g3768 ( .o(n9256), .a(n8178) );
in01f01  g3769 ( .o(n9257), .a(n8179) );
na02f01  g3770 ( .o(n9258), .a(n9257), .b(n8160_1) );
na02f01  g3771 ( .o(n9259), .a(n9258), .b(n9256) );
no02f01  g3772 ( .o(n9260), .a(n9259), .b(n9255) );
no02f01  g3773 ( .o(n9261), .a(n5719_1), .b(n7005) );
no02f01  g3774 ( .o(n9262), .a(_net_9933), .b(_net_10369) );
no02f01  g3775 ( .o(n9263), .a(n9262), .b(n9261) );
in01f01  g3776 ( .o(n9264), .a(n9263) );
ao12f01  g3777 ( .o(n9265), .a(n8184), .b(n9264), .c(n9260) );
oa12f01  g3778 ( .o(n9266), .a(n9265), .b(n9264), .c(n9260) );
no02f01  g3779 ( .o(n9267), .a(n8196), .b(_net_10369) );
in01f01  g3780 ( .o(n9268), .a(n9267) );
na02f01  g3781 ( .o(n9269), .a(n8196), .b(_net_10369) );
na02f01  g3782 ( .o(n9270), .a(n9269), .b(n9268) );
ao22f01  g3783 ( .o(n9271), .a(n9270), .b(n8200_1), .c(n8202), .d(_net_10369) );
na02f01  g3784 ( .o(n1965), .a(n9271), .b(n9266) );
na02f01  g3785 ( .o(n9273), .a(n7358), .b(net_253) );
na02f01  g3786 ( .o(n9274), .a(n7352), .b(net_9684) );
ao22f01  g3787 ( .o(n9275), .a(n7357), .b(_net_10117), .c(n7353), .d(x4587) );
na04f01  g3788 ( .o(n1970), .a(n9275), .b(n9274), .c(n9273), .d(n7355_1) );
in01f01  g3789 ( .o(n9277), .a(n6632) );
no02f01  g3790 ( .o(n9278), .a(n6640), .b(n6618) );
in01f01  g3791 ( .o(n9279), .a(n9278) );
na02f01  g3792 ( .o(n9280), .a(n9279), .b(n9277) );
na02f01  g3793 ( .o(n9281), .a(n9278), .b(n6632) );
na02f01  g3794 ( .o(n1975), .a(n9281), .b(n9280) );
no02f01  g3795 ( .o(n1980), .a(net_9613), .b(net_9614) );
na02f01  g3796 ( .o(n9284), .a(net_9348), .b(n7890) );
in01f01  g3797 ( .o(n9285), .a(net_9348) );
na02f01  g3798 ( .o(n9286), .a(n9285), .b(_net_9344) );
na02f01  g3799 ( .o(n9287), .a(n6454), .b(net_9347) );
in01f01  g3800 ( .o(n9288), .a(net_9347) );
na02f01  g3801 ( .o(n9289), .a(_net_9343), .b(n9288) );
ao22f01  g3802 ( .o(n9290), .a(n9289), .b(n9287), .c(n9286), .d(n9284) );
na02f01  g3803 ( .o(n9291), .a(net_9349), .b(n6457) );
in01f01  g3804 ( .o(n9292), .a(net_9349) );
na02f01  g3805 ( .o(n9293), .a(n9292), .b(_net_9345) );
na02f01  g3806 ( .o(n9294), .a(net_9350), .b(n7730) );
in01f01  g3807 ( .o(n9295), .a(net_9350) );
na02f01  g3808 ( .o(n9296), .a(n9295), .b(_net_9346) );
ao22f01  g3809 ( .o(n9297), .a(n9296), .b(n9294), .c(n9293), .d(n9291) );
na02f01  g3810 ( .o(n1985), .a(n9297), .b(n9290) );
na02f01  g3811 ( .o(n9299), .a(n6038), .b(net_262) );
na02f01  g3812 ( .o(n9300), .a(n6037_1), .b(net_9891) );
ao22f01  g3813 ( .o(n9301), .a(n6044), .b(x3889), .c(n6042_1), .d(_net_10336) );
na04f01  g3814 ( .o(n1990), .a(n9301), .b(n9300), .c(n9299), .d(n6040) );
ao12f01  g3815 ( .o(n9303), .a(n5658), .b(n6532), .c(net_238) );
ao22f01  g3816 ( .o(n9304), .a(n6535), .b(x5647), .c(n6534), .d(net_9998) );
na02f01  g3817 ( .o(n1995), .a(n9304), .b(n9303) );
na03f01  g3818 ( .o(n9306), .a(n7663), .b(n8219_1), .c(n7361) );
na04f01  g3819 ( .o(n9307), .a(n9044), .b(n9041), .c(n9043), .d(n8793) );
no04f01  g3820 ( .o(n9308), .a(n9307), .b(n9306), .c(_net_10436), .d(_net_10435) );
no03f01  g3821 ( .o(n2000), .a(n9308), .b(_net_10049), .c(n9055) );
ao12f01  g3822 ( .o(n9310), .a(n5658), .b(n7844), .c(net_246) );
ao22f01  g3823 ( .o(n9311), .a(n7847), .b(x5143), .c(n7846), .d(net_9808) );
na02f01  g3824 ( .o(n2005), .a(n9311), .b(n9310) );
ao12f01  g3825 ( .o(n9313), .a(n5658), .b(n6532), .c(net_236) );
ao22f01  g3826 ( .o(n9314), .a(n6535), .b(x5790), .c(n6534), .d(net_9996) );
na02f01  g3827 ( .o(n2010), .a(n9314), .b(n9313) );
no02f01  g3828 ( .o(n9316), .a(n7678), .b(_net_10439) );
na02f01  g3829 ( .o(n9317), .a(n9316), .b(n8793) );
in01f01  g3830 ( .o(n9318), .a(n9316) );
na02f01  g3831 ( .o(n9319), .a(n9318), .b(_net_10440) );
na02f01  g3832 ( .o(n2015), .a(n9319), .b(n9317) );
in01f01  g3833 ( .o(n9321), .a(_net_10373) );
no02f01  g3834 ( .o(n9322), .a(n5705_1), .b(n7003_1) );
no02f01  g3835 ( .o(n9323), .a(_net_9934), .b(_net_10370) );
in01f01  g3836 ( .o(n9324), .a(n9323) );
na02f01  g3837 ( .o(n9325), .a(n5719_1), .b(n7005) );
oa12f01  g3838 ( .o(n9326), .a(n9325), .b(n9261), .c(n8178) );
na02f01  g3839 ( .o(n9327), .a(n9326), .b(n9258) );
no02f01  g3840 ( .o(n9328), .a(n9327), .b(n9255) );
oa22f01  g3841 ( .o(n9329), .a(n9328), .b(n9262), .c(n9326), .d(n7005) );
ao12f01  g3842 ( .o(n9330), .a(n9322), .b(n9329), .c(n9324) );
no02f01  g3843 ( .o(n9331), .a(n9330), .b(n6996) );
na02f01  g3844 ( .o(n9332), .a(n9331), .b(_net_10372) );
ao12f01  g3845 ( .o(n9333), .a(n8184), .b(n9332), .c(n9321) );
oa12f01  g3846 ( .o(n9334), .a(n9333), .b(n9332), .c(n9321) );
na02f01  g3847 ( .o(n9335), .a(n9267), .b(n7003_1) );
no02f01  g3848 ( .o(n9336), .a(n9335), .b(_net_10371) );
na03f01  g3849 ( .o(n9337), .a(n9336), .b(n7062), .c(_net_10373) );
ao12f01  g3850 ( .o(n9338), .a(_net_10373), .b(n9336), .c(n7062) );
no02f01  g3851 ( .o(n9339), .a(n9338), .b(n9144) );
ao22f01  g3852 ( .o(n9340), .a(n9339), .b(n9337), .c(n8202), .d(_net_10373) );
na02f01  g3853 ( .o(n2020), .a(n9340), .b(n9334) );
no03f01  g3854 ( .o(n9342), .a(n6812), .b(n6810), .c(n6803) );
no02f01  g3855 ( .o(n9343), .a(n6814), .b(n6777) );
in01f01  g3856 ( .o(n9344), .a(n9343) );
ao12f01  g3857 ( .o(n9345), .a(n6933), .b(n9344), .c(n9342) );
oa12f01  g3858 ( .o(n9346), .a(n9345), .b(n9344), .c(n9342) );
na02f01  g3859 ( .o(n9347), .a(n6839), .b(n6813) );
no02f01  g3860 ( .o(n9348), .a(n6840), .b(n6846_1) );
ao22f01  g3861 ( .o(n9349), .a(n9348), .b(n9347), .c(n6168), .d(_net_10252) );
na02f01  g3862 ( .o(n2025), .a(n9349), .b(n9346) );
in01f01  g3863 ( .o(n9351), .a(net_10290) );
no02f01  g3864 ( .o(n9352), .a(n7464), .b(n6884) );
na02f01  g3865 ( .o(n9353), .a(n7466), .b(n6883) );
oa22f01  g3866 ( .o(n2030), .a(n9353), .b(n5546), .c(n9352), .d(n9351) );
na03f01  g3867 ( .o(n9355), .a(_net_10430), .b(_net_10431), .c(_net_10429) );
na02f01  g3868 ( .o(n2035), .a(n9355), .b(n7666) );
in01f01  g3869 ( .o(n9357), .a(n7821_1) );
ao12f01  g3870 ( .o(n9358), .a(n7823), .b(n9357), .c(n7762) );
in01f01  g3871 ( .o(n9359), .a(n9358) );
ao12f01  g3872 ( .o(n9360), .a(n9359), .b(n9357), .c(n7818) );
in01f01  g3873 ( .o(n9361), .a(_net_10162) );
no02f01  g3874 ( .o(n9362), .a(n9361), .b(_net_10124) );
in01f01  g3875 ( .o(n9363), .a(_net_10124) );
no02f01  g3876 ( .o(n9364), .a(_net_10162), .b(n9363) );
no02f01  g3877 ( .o(n9365), .a(n9364), .b(n9362) );
na02f01  g3878 ( .o(n9366), .a(n9365), .b(n9360) );
in01f01  g3879 ( .o(n9367), .a(n9360) );
in01f01  g3880 ( .o(n9368), .a(n9365) );
na02f01  g3881 ( .o(n9369), .a(n9368), .b(n9367) );
na02f01  g3882 ( .o(n2040), .a(n9369), .b(n9366) );
no02f01  g3883 ( .o(n9371), .a(n8762_1), .b(_net_9325) );
no02f01  g3884 ( .o(n9372), .a(_net_9324), .b(n7882) );
no02f01  g3885 ( .o(n9373), .a(n9372), .b(n9371) );
no02f01  g3886 ( .o(n9374), .a(net_9153), .b(n8984) );
in01f01  g3887 ( .o(n9375), .a(net_9153) );
no02f01  g3888 ( .o(n9376), .a(n9375), .b(net_9154) );
no02f01  g3889 ( .o(n9377), .a(n9376), .b(n9374) );
na02f01  g3890 ( .o(n9378), .a(n9377), .b(n9373) );
in01f01  g3891 ( .o(n9379), .a(n9373) );
in01f01  g3892 ( .o(n9380), .a(n9377) );
na02f01  g3893 ( .o(n9381), .a(n9380), .b(n9379) );
na03f01  g3894 ( .o(n9382), .a(n9381), .b(n9378), .c(n8638) );
ao12f01  g3895 ( .o(n9383), .a(n7883), .b(n8637), .c(_net_9318) );
na02f01  g3896 ( .o(n2045), .a(n9383), .b(n9382) );
in01f01  g3897 ( .o(n9385), .a(_net_9850) );
oa22f01  g3898 ( .o(n2050), .a(n7480_1), .b(n9385), .c(n7478), .d(n5609) );
ao12f01  g3899 ( .o(n9387), .a(n5658), .b(n6875_1), .c(net_240) );
ao22f01  g3900 ( .o(n9388), .a(n6878), .b(x5548), .c(n6877), .d(net_9901) );
na02f01  g3901 ( .o(n2055), .a(n9388), .b(n9387) );
na02f01  g3902 ( .o(n9390), .a(n7958), .b(_net_8828) );
ao12f01  g3903 ( .o(n2060), .a(n5658), .b(n9390), .c(n8746) );
no02f01  g3904 ( .o(n9392), .a(n8267), .b(_net_202) );
na02f01  g3905 ( .o(n9393), .a(n8270), .b(n573) );
oa22f01  g3906 ( .o(n2065), .a(n9393), .b(n9392), .c(n8280), .d(n8258) );
in01f01  g3907 ( .o(n9395), .a(_net_9213) );
no02f01  g3908 ( .o(n9396), .a(n6686), .b(net_9218) );
na02f01  g3909 ( .o(n9397), .a(n9396), .b(net_9227) );
no02f01  g3910 ( .o(n9398), .a(n8091_1), .b(n8547) );
in01f01  g3911 ( .o(n9399), .a(n9398) );
no02f01  g3912 ( .o(n9400), .a(n9399), .b(n8090) );
in01f01  g3913 ( .o(n9401), .a(n9400) );
na02f01  g3914 ( .o(n9402), .a(n9401), .b(n9395) );
no02f01  g3915 ( .o(n9403), .a(n9401), .b(n9395) );
in01f01  g3916 ( .o(n9404), .a(n9403) );
na02f01  g3917 ( .o(n9405), .a(n9404), .b(n9402) );
in01f01  g3918 ( .o(n9406), .a(net_9227) );
na02f01  g3919 ( .o(n9407), .a(n9396), .b(n9406) );
oa22f01  g3920 ( .o(n2075), .a(n9407), .b(n9395), .c(n9405), .d(n9397) );
in01f01  g3921 ( .o(n9409), .a(net_9511) );
ao22f01  g3922 ( .o(n9410), .a(n8118), .b(x2826), .c(n8117), .d(_net_9396) );
oa12f01  g3923 ( .o(n2080), .a(n9410), .b(n8116_1), .c(n9409) );
na04f01  g3924 ( .o(n9412), .a(n6570), .b(n6558), .c(n5663), .d(x6496) );
in01f01  g3925 ( .o(n9413), .a(_net_8847) );
na02f01  g3926 ( .o(n9414), .a(n9413), .b(_net_10528) );
ao12f01  g3927 ( .o(n2085), .a(n5658), .b(n9414), .c(n9412) );
na02f01  g3928 ( .o(n9416), .a(net_106), .b(net_107) );
na02f01  g3929 ( .o(n9417), .a(net_101), .b(net_103) );
no02f01  g3930 ( .o(n9418), .a(n9417), .b(n9416) );
na03f01  g3931 ( .o(n9419), .a(n9418), .b(net_100), .c(net_116) );
na04f01  g3932 ( .o(n9420), .a(net_105), .b(net_110), .c(net_102), .d(net_111) );
na04f01  g3933 ( .o(n9421), .a(net_113), .b(net_114), .c(net_104), .d(net_109) );
no02f01  g3934 ( .o(n9422), .a(n9421), .b(n9420) );
na04f01  g3935 ( .o(n9423), .a(n9422), .b(net_108), .c(net_112), .d(net_115) );
no02f01  g3936 ( .o(n2090), .a(n9423), .b(n9419) );
ao12f01  g3937 ( .o(n9425), .a(n5658), .b(n6887), .c(x4449) );
oa12f01  g3938 ( .o(n2095), .a(n9425), .b(n6885_1), .c(n9198) );
ao12f01  g3939 ( .o(n9427), .a(n5658), .b(n6160_1), .c(x4117) );
oa12f01  g3940 ( .o(n2100), .a(n9427), .b(n6159), .c(n7822) );
ao12f01  g3941 ( .o(n9429), .a(n5658), .b(n6052_1), .c(x4359) );
oa12f01  g3942 ( .o(n2105), .a(n9429), .b(n6048), .c(n8240_1) );
in01f01  g3943 ( .o(n9431), .a(_net_10103) );
ao12f01  g3944 ( .o(n9432), .a(n5658), .b(n6160_1), .c(x5601) );
oa12f01  g3945 ( .o(n2110), .a(n9432), .b(n6159), .c(n9431) );
in01f01  g3946 ( .o(n9434), .a(_net_10098) );
ao12f01  g3947 ( .o(n9435), .a(n5658), .b(n6160_1), .c(x5901) );
oa12f01  g3948 ( .o(n2115), .a(n9435), .b(n6159), .c(n9434) );
no02f01  g3949 ( .o(n9437), .a(n6910_1), .b(n6909) );
no02f01  g3950 ( .o(n9438), .a(n9437), .b(n6919_1) );
no02f01  g3951 ( .o(n9439), .a(n6917), .b(n6912) );
in01f01  g3952 ( .o(n9440), .a(n9439) );
ao12f01  g3953 ( .o(n9441), .a(n6933), .b(n9440), .c(n9438) );
oa12f01  g3954 ( .o(n9442), .a(n9441), .b(n9440), .c(n9438) );
na02f01  g3955 ( .o(n9443), .a(n6940), .b(_net_10262) );
na02f01  g3956 ( .o(n9444), .a(n9443), .b(n6942) );
ao22f01  g3957 ( .o(n9445), .a(n9444), .b(n6175), .c(n6168), .d(_net_10262) );
na02f01  g3958 ( .o(n2120), .a(n9445), .b(n9442) );
in01f01  g3959 ( .o(n9447), .a(net_208) );
in01f01  g3960 ( .o(n9448), .a(net_207) );
no02f01  g3961 ( .o(n9449), .a(n8276_1), .b(n9448) );
in01f01  g3962 ( .o(n9450), .a(n9449) );
no02f01  g3963 ( .o(n9451), .a(n9450), .b(n9447) );
oa12f01  g3964 ( .o(n9452), .a(n573), .b(n9449), .c(net_208) );
oa22f01  g3965 ( .o(n2125), .a(n9452), .b(n9451), .c(n8280), .d(n9447) );
in01f01  g3966 ( .o(n9454), .a(n7991) );
in01f01  g3967 ( .o(n9455), .a(net_9527) );
in01f01  g3968 ( .o(n9456), .a(net_9525) );
in01f01  g3969 ( .o(n9457), .a(net_9524) );
in01f01  g3970 ( .o(n9458), .a(net_9522) );
in01f01  g3971 ( .o(n9459), .a(_net_9520) );
no02f01  g3972 ( .o(n9460), .a(n7996_1), .b(_net_9519) );
na02f01  g3973 ( .o(n9461), .a(n9460), .b(n9459) );
no02f01  g3974 ( .o(n9462), .a(n9461), .b(_net_9521) );
na02f01  g3975 ( .o(n9463), .a(n9462), .b(n9458) );
no02f01  g3976 ( .o(n9464), .a(n9463), .b(net_9523) );
na03f01  g3977 ( .o(n9465), .a(n9464), .b(n9457), .c(n9456) );
no02f01  g3978 ( .o(n9466), .a(n9465), .b(net_9526) );
na02f01  g3979 ( .o(n9467), .a(n9466), .b(n9455) );
no02f01  g3980 ( .o(n9468), .a(n9467), .b(net_9528) );
in01f01  g3981 ( .o(n9469), .a(n9468) );
na02f01  g3982 ( .o(n9470), .a(n9467), .b(net_9528) );
ao12f01  g3983 ( .o(n9471), .a(n7999), .b(n9470), .c(n9469) );
in01f01  g3984 ( .o(n9472), .a(net_9528) );
oa12f01  g3985 ( .o(n9473), .a(x6599), .b(n8002), .c(n9472) );
no02f01  g3986 ( .o(n9474), .a(n9473), .b(n9471) );
oa12f01  g3987 ( .o(n2135), .a(n9474), .b(n8929), .c(n9454) );
na02f01  g3988 ( .o(n9476), .a(n7937), .b(_net_231) );
na02f01  g3989 ( .o(n9477), .a(n7936), .b(net_9761) );
ao22f01  g3990 ( .o(n9478), .a(n7943), .b(_net_10200), .c(n7942), .d(x6102) );
na04f01  g3991 ( .o(n2145), .a(n9478), .b(n9477), .c(n9476), .d(n7939) );
na02f01  g3992 ( .o(n9480), .a(n6056), .b(net_244) );
na02f01  g3993 ( .o(n9481), .a(n6055), .b(net_9972) );
ao22f01  g3994 ( .o(n9482), .a(n6062_1), .b(x5289), .c(n6060), .d(_net_10423) );
na04f01  g3995 ( .o(n2150), .a(n9482), .b(n9481), .c(n9480), .d(n6058) );
ao12f01  g3996 ( .o(n9484), .a(n5658), .b(n6875_1), .c(_net_233) );
ao22f01  g3997 ( .o(n9485), .a(n6878), .b(x5961), .c(n6877), .d(net_9894) );
na02f01  g3998 ( .o(n2155), .a(n9485), .b(n9484) );
ao12f01  g3999 ( .o(n9487), .a(n7975), .b(n8748), .c(_net_9639) );
no04f01  g4000 ( .o(n9488), .a(n9487), .b(n8751), .c(n7969), .d(n7964) );
in01f01  g4001 ( .o(n9489), .a(_net_9639) );
in01f01  g4002 ( .o(n9490), .a(n8769) );
no04f01  g4003 ( .o(n9491), .a(n9490), .b(n8752), .c(n8753), .d(n9489) );
in01f01  g4004 ( .o(n9492), .a(net_9612) );
na04f01  g4005 ( .o(n9493), .a(n8774), .b(n9492), .c(_net_9640), .d(_net_9639) );
in01f01  g4006 ( .o(n9494), .a(n7972_1) );
no02f01  g4007 ( .o(n9495), .a(n9494), .b(n8744) );
no02f01  g4008 ( .o(n9496), .a(net_9279), .b(n9489) );
no02f01  g4009 ( .o(n9497), .a(n9496), .b(n9495) );
oa12f01  g4010 ( .o(n9498), .a(n9493), .b(n9497), .c(n9489) );
no03f01  g4011 ( .o(n9499), .a(n9498), .b(n9491), .c(n9488) );
na02f01  g4012 ( .o(n9500), .a(n8743), .b(x6599) );
no02f01  g4013 ( .o(n2165), .a(n9500), .b(n9499) );
in01f01  g4014 ( .o(n9502), .a(n8214_1) );
na02f01  g4015 ( .o(n9503), .a(n8236), .b(n9502) );
no02f01  g4016 ( .o(n9504), .a(n8211), .b(n8210_1) );
in01f01  g4017 ( .o(n9505), .a(n9504) );
na02f01  g4018 ( .o(n9506), .a(n9505), .b(n9503) );
na03f01  g4019 ( .o(n9507), .a(n9504), .b(n8236), .c(n9502) );
na02f01  g4020 ( .o(n2174), .a(n9507), .b(n9506) );
ao12f01  g4021 ( .o(n9509), .a(n5658), .b(n6875_1), .c(net_252) );
ao22f01  g4022 ( .o(n9510), .a(n6878), .b(x4694), .c(n6877), .d(net_9913) );
na02f01  g4023 ( .o(n2179), .a(n9510), .b(n9509) );
ao22f01  g4024 ( .o(n9512), .a(n5842), .b(net_9687), .c(n5841), .d(_net_125) );
na02f01  g4025 ( .o(n9513), .a(n5847), .b(net_9984) );
ao22f01  g4026 ( .o(n9514), .a(n5850), .b(net_9786), .c(n5849_1), .d(net_9885) );
na03f01  g4027 ( .o(n2184), .a(n9514), .b(n9513), .c(n9512) );
in01f01  g4028 ( .o(n9516), .a(net_10039) );
oa22f01  g4029 ( .o(n2193), .a(n5907), .b(n9516), .c(n5905), .d(n5591) );
in01f01  g4030 ( .o(n9518), .a(net_214) );
oa22f01  g4031 ( .o(n2198), .a(n7756), .b(n6407), .c(n7755), .d(n9518) );
no02f01  g4032 ( .o(n9520), .a(n6632), .b(n6618) );
no02f01  g4033 ( .o(n9521), .a(n6639_1), .b(n6637) );
in01f01  g4034 ( .o(n9522), .a(n9521) );
oa12f01  g4035 ( .o(n9523), .a(n9522), .b(n6640), .c(n9520) );
in01f01  g4036 ( .o(n9524), .a(n9520) );
in01f01  g4037 ( .o(n9525), .a(n6640) );
na03f01  g4038 ( .o(n9526), .a(n9521), .b(n9525), .c(n9524) );
na02f01  g4039 ( .o(n2207), .a(n9526), .b(n9523) );
in01f01  g4040 ( .o(n9528), .a(_net_10311) );
ao12f01  g4041 ( .o(n9529), .a(n5658), .b(n5774), .c(x5722) );
oa12f01  g4042 ( .o(n2212), .a(n9529), .b(n5770), .c(n9528) );
in01f01  g4043 ( .o(n9531), .a(net_10050) );
oa12f01  g4044 ( .o(n9532), .a(x6599), .b(n8828), .c(n6529) );
na02f01  g4045 ( .o(n9533), .a(n8830), .b(net_10490) );
oa22f01  g4046 ( .o(n2222), .a(n9533), .b(n8827), .c(n9532), .d(n9531) );
in01f01  g4047 ( .o(n9535), .a(_net_10413) );
ao12f01  g4048 ( .o(n9536), .a(n5658), .b(n6052_1), .c(x5901) );
oa12f01  g4049 ( .o(n2232), .a(n9536), .b(n6048), .c(n9535) );
oa22f01  g4050 ( .o(n2237), .a(n7756), .b(n6387), .c(n7755), .d(n8284) );
in01f01  g4051 ( .o(n9539), .a(n8749) );
na02f01  g4052 ( .o(n9540), .a(n8750), .b(n9539) );
no03f01  g4053 ( .o(n9541), .a(n9540), .b(n7966), .c(n8772_1) );
no02f01  g4054 ( .o(n9542), .a(n9490), .b(n8752) );
na03f01  g4055 ( .o(n9543), .a(n9542), .b(_net_9641), .c(_net_9640) );
in01f01  g4056 ( .o(n9544), .a(n9497) );
no02f01  g4057 ( .o(n9545), .a(net_9612), .b(n8772_1) );
in01f01  g4058 ( .o(n9546), .a(n9545) );
no02f01  g4059 ( .o(n9547), .a(n9546), .b(n8773) );
oa12f01  g4060 ( .o(n9548), .a(_net_9640), .b(n9547), .c(n9544) );
in01f01  g4061 ( .o(n9549), .a(_net_185) );
no02f01  g4062 ( .o(n9550), .a(net_186), .b(n9549) );
in01f01  g4063 ( .o(n9551), .a(n9550) );
na03f01  g4064 ( .o(n9552), .a(n9551), .b(net_9279), .c(_net_9639) );
na03f01  g4065 ( .o(n9553), .a(n9552), .b(n9548), .c(n9543) );
oa12f01  g4066 ( .o(n9554), .a(x6599), .b(n9553), .c(n9541) );
no02f01  g4067 ( .o(n2242), .a(n9554), .b(n2827) );
no03f01  g4068 ( .o(n9556), .a(n9111), .b(n9109), .c(n9103) );
in01f01  g4069 ( .o(n9557), .a(n9556) );
no02f01  g4070 ( .o(n9558), .a(n9113), .b(n9082) );
ao12f01  g4071 ( .o(n9559), .a(n8184), .b(n9558), .c(n9557) );
oa12f01  g4072 ( .o(n9560), .a(n9559), .b(n9558), .c(n9557) );
na02f01  g4073 ( .o(n9561), .a(n9139), .b(n9112) );
no02f01  g4074 ( .o(n9562), .a(n9140), .b(n9144) );
ao22f01  g4075 ( .o(n9563), .a(n9562), .b(n9561), .c(n8202), .d(_net_10357) );
na02f01  g4076 ( .o(n2251), .a(n9563), .b(n9560) );
no02f01  g4077 ( .o(n2690), .a(n6021), .b(n8897) );
in01f01  g4078 ( .o(n9566), .a(n2690) );
in01f01  g4079 ( .o(n9567), .a(n9466) );
na02f01  g4080 ( .o(n9568), .a(n9567), .b(net_9527) );
ao12f01  g4081 ( .o(n9569), .a(n7999), .b(n9568), .c(n9467) );
oa12f01  g4082 ( .o(n9570), .a(x6599), .b(n8002), .c(n9455) );
no02f01  g4083 ( .o(n9571), .a(n9570), .b(n9569) );
oa12f01  g4084 ( .o(n2256), .a(n9571), .b(n9566), .c(n9454) );
na02f01  g4085 ( .o(n9573), .a(n6038), .b(net_249) );
na02f01  g4086 ( .o(n9574), .a(n6037_1), .b(net_9878) );
ao22f01  g4087 ( .o(n9575), .a(n6044), .b(x4937), .c(n6042_1), .d(_net_10323) );
na04f01  g4088 ( .o(n2261), .a(n9575), .b(n9574), .c(n9573), .d(n6040) );
in01f01  g4089 ( .o(n9577), .a(net_215) );
oa22f01  g4090 ( .o(n2266), .a(n7756), .b(n6373_1), .c(n7755), .d(n9577) );
in01f01  g4091 ( .o(n9579), .a(_net_9949) );
na03f01  g4092 ( .o(n9580), .a(n8932), .b(n7017_1), .c(n7018) );
na04f01  g4093 ( .o(n9581), .a(n6999), .b(n7064), .c(n6994), .d(n8931) );
no04f01  g4094 ( .o(n9582), .a(n9581), .b(n9580), .c(_net_10330), .d(_net_10331) );
no03f01  g4095 ( .o(n2271), .a(n9582), .b(_net_9950), .c(n9579) );
ao12f01  g4096 ( .o(n9584), .a(n5658), .b(n6887), .c(x4285) );
oa12f01  g4097 ( .o(n2276), .a(n9584), .b(n6885_1), .c(n9204) );
na02f01  g4098 ( .o(n9586), .a(n6056), .b(_net_234) );
na02f01  g4099 ( .o(n9587), .a(n6055), .b(net_9962) );
ao22f01  g4100 ( .o(n9588), .a(n6062_1), .b(x5901), .c(n6060), .d(_net_10413) );
na04f01  g4101 ( .o(n2281), .a(n9588), .b(n9587), .c(n9586), .d(n6058) );
na02f01  g4102 ( .o(n9590), .a(n6038), .b(_net_254) );
na02f01  g4103 ( .o(n9591), .a(n6037_1), .b(net_9883) );
ao22f01  g4104 ( .o(n9592), .a(n6044), .b(x4520), .c(n6042_1), .d(_net_10328) );
na04f01  g4105 ( .o(n2286), .a(n9592), .b(n9591), .c(n9590), .d(n6040) );
na03f01  g4106 ( .o(n9594), .a(_net_9503), .b(n8399_1), .c(net_9533) );
oa12f01  g4107 ( .o(n9595), .a(n5738), .b(_net_8955), .c(_net_9062) );
ao12f01  g4108 ( .o(n2291), .a(n9595), .b(n9594), .c(n5884) );
ao12f01  g4109 ( .o(n9597), .a(n5658), .b(n5678), .c(net_247) );
ao22f01  g4110 ( .o(n9598), .a(n5681_1), .b(x5077), .c(n5680), .d(net_9710) );
na02f01  g4111 ( .o(n2296), .a(n9598), .b(n9597) );
in01f01  g4112 ( .o(n9600), .a(net_10194) );
na02f01  g4113 ( .o(n9601), .a(net_263), .b(net_10175) );
ao12f01  g4114 ( .o(n2301), .a(n8577_1), .b(n9601), .c(n9600) );
in01f01  g4115 ( .o(n9603), .a(n8704) );
no02f01  g4116 ( .o(n9604), .a(n9603), .b(net_9653) );
no03f01  g4117 ( .o(n2306), .a(n9604), .b(n8706), .c(net_9151) );
na02f01  g4118 ( .o(n9606), .a(n7453), .b(_net_10468) );
no02f01  g4119 ( .o(n9607), .a(n7395), .b(n7398_1) );
oa12f01  g4120 ( .o(n9608), .a(n7450), .b(n9607), .c(n7434) );
in01f01  g4121 ( .o(n9609), .a(n7397) );
na03f01  g4122 ( .o(n9610), .a(n7402), .b(n7400), .c(n9609) );
oa12f01  g4123 ( .o(n9611), .a(n8066), .b(n7401), .c(n7397) );
na03f01  g4124 ( .o(n9612), .a(n9611), .b(n9610), .c(n7431) );
na03f01  g4125 ( .o(n2311), .a(n9612), .b(n9608), .c(n9606) );
ao12f01  g4126 ( .o(n9614), .a(n5658), .b(n7844), .c(_net_232) );
ao22f01  g4127 ( .o(n9615), .a(n7847), .b(x6028), .c(n7846), .d(net_9794) );
na02f01  g4128 ( .o(n2316), .a(n9615), .b(n9614) );
na02f01  g4129 ( .o(n9617), .a(n6020), .b(n5994) );
oa12f01  g4130 ( .o(n7418), .a(n9617), .b(n6020), .c(n5990) );
na02f01  g4131 ( .o(n9619), .a(n7418), .b(n7991) );
in01f01  g4132 ( .o(n9620), .a(n9464) );
no03f01  g4133 ( .o(n9621), .a(n9620), .b(net_9524), .c(net_9525) );
ao12f01  g4134 ( .o(n9622), .a(n9456), .b(n9464), .c(n9457) );
oa12f01  g4135 ( .o(n9623), .a(n7998), .b(n9622), .c(n9621) );
no02f01  g4136 ( .o(n9624), .a(n8002), .b(n9456) );
no02f01  g4137 ( .o(n9625), .a(n9624), .b(n5658) );
na03f01  g4138 ( .o(n2321), .a(n9625), .b(n9623), .c(n9619) );
no03f01  g4139 ( .o(n2330), .a(n2827), .b(n7915), .c(n6354) );
ao22f01  g4140 ( .o(n9628), .a(n5842), .b(net_9709), .c(n5841), .d(net_149) );
na02f01  g4141 ( .o(n9629), .a(n5847), .b(net_10006) );
ao22f01  g4142 ( .o(n9630), .a(n5850), .b(net_9808), .c(n5849_1), .d(net_9907) );
na03f01  g4143 ( .o(n2342), .a(n9630), .b(n9629), .c(n9628) );
in01f01  g4144 ( .o(n9632), .a(x3638) );
no02f01  g4145 ( .o(n2347), .a(n9632), .b(n5658) );
in01f01  g4146 ( .o(n9634), .a(n9330) );
no02f01  g4147 ( .o(n9635), .a(n9634), .b(n6996) );
no02f01  g4148 ( .o(n9636), .a(n9330), .b(_net_10371) );
oa12f01  g4149 ( .o(n9637), .a(n8183), .b(n9636), .c(n9635) );
no02f01  g4150 ( .o(n9638), .a(n9335), .b(n6996) );
ao12f01  g4151 ( .o(n9639), .a(_net_10371), .b(n9267), .c(n7003_1) );
no03f01  g4152 ( .o(n9640), .a(n9639), .b(n9638), .c(n9144) );
ao12f01  g4153 ( .o(n9641), .a(n9640), .b(n8202), .c(_net_10371) );
na02f01  g4154 ( .o(n2352), .a(n9641), .b(n9637) );
na02f01  g4155 ( .o(n9643), .a(n7358), .b(net_248) );
na02f01  g4156 ( .o(n9644), .a(n7352), .b(net_9679) );
ao22f01  g4157 ( .o(n9645), .a(n7357), .b(_net_10112), .c(n7353), .d(x5003) );
na04f01  g4158 ( .o(n2357), .a(n9645), .b(n9644), .c(n9643), .d(n7355_1) );
ao12f01  g4159 ( .o(n9647), .a(n5658), .b(n6875_1), .c(net_239) );
ao22f01  g4160 ( .o(n9648), .a(n6878), .b(x5601), .c(n6877), .d(net_9900) );
na02f01  g4161 ( .o(n2362), .a(n9648), .b(n9647) );
ao22f01  g4162 ( .o(n9650), .a(n5842), .b(net_9692), .c(n5841), .d(_net_130) );
na02f01  g4163 ( .o(n9651), .a(n5847), .b(net_9989) );
ao22f01  g4164 ( .o(n9652), .a(n5850), .b(net_9791), .c(n5849_1), .d(net_9890) );
na03f01  g4165 ( .o(n2375), .a(n9652), .b(n9651), .c(n9650) );
oa22f01  g4166 ( .o(n2380), .a(n5694), .b(n8181), .c(n5692), .d(n5582_1) );
in01f01  g4167 ( .o(n9655), .a(_net_9752) );
no02f01  g4168 ( .o(n9656), .a(n9655), .b(_net_9751) );
in01f01  g4169 ( .o(n9657), .a(n9656) );
in01f01  g4170 ( .o(n9658), .a(_net_10163) );
no03f01  g4171 ( .o(n9659), .a(_net_10162), .b(_net_10160), .c(_net_10155) );
na03f01  g4172 ( .o(n9660), .a(n9659), .b(n7820), .c(n9658) );
no04f01  g4173 ( .o(n9661), .a(_net_10157), .b(_net_10159), .c(_net_10158), .d(_net_10156) );
na02f01  g4174 ( .o(n9662), .a(n9661), .b(n7778_1) );
no02f01  g4175 ( .o(n9663), .a(n9662), .b(n9660) );
no02f01  g4176 ( .o(n2385), .a(n9663), .b(n9657) );
in01f01  g4177 ( .o(n9665), .a(net_10508) );
in01f01  g4178 ( .o(n9666), .a(net_10503) );
na02f01  g4179 ( .o(n9667), .a(n9666), .b(x6599) );
na02f01  g4180 ( .o(n9668), .a(n8580), .b(net_10490) );
ao12f01  g4181 ( .o(n2390), .a(n9667), .b(n9668), .c(n9665) );
no02f01  g4182 ( .o(n9670), .a(n5986), .b(net_9598) );
in01f01  g4183 ( .o(n9671), .a(n9670) );
in01f01  g4184 ( .o(n9672), .a(n6658) );
ao12f01  g4185 ( .o(n9673), .a(n6659_1), .b(n9672), .c(n6611) );
in01f01  g4186 ( .o(n9674), .a(n9673) );
in01f01  g4187 ( .o(n9675), .a(n6615) );
oa12f01  g4188 ( .o(n9676), .a(n9675), .b(n6648), .c(n6638) );
no02f01  g4189 ( .o(n9677), .a(n6658), .b(n6655) );
in01f01  g4190 ( .o(n9678), .a(n9677) );
ao12f01  g4191 ( .o(n9679), .a(n9678), .b(n6651), .c(n9676) );
na02f01  g4192 ( .o(n9680), .a(n5986), .b(net_9598) );
oa12f01  g4193 ( .o(n9681), .a(n9680), .b(n9679), .c(n9674) );
na02f01  g4194 ( .o(n9682), .a(n9681), .b(n9671) );
in01f01  g4195 ( .o(n9683), .a(net_9599) );
no02f01  g4196 ( .o(n9684), .a(n6011), .b(n9683) );
no02f01  g4197 ( .o(n9685), .a(n8897), .b(net_9599) );
no02f01  g4198 ( .o(n9686), .a(n9685), .b(n9684) );
in01f01  g4199 ( .o(n9687), .a(n9686) );
na02f01  g4200 ( .o(n9688), .a(n9687), .b(n9682) );
na03f01  g4201 ( .o(n9689), .a(n9686), .b(n9681), .c(n9671) );
na02f01  g4202 ( .o(n2395), .a(n9689), .b(n9688) );
in01f01  g4203 ( .o(n9691), .a(net_9750) );
oa22f01  g4204 ( .o(n2400), .a(n7367), .b(n9691), .c(n7365_1), .d(n5567_1) );
na02f01  g4205 ( .o(n9693), .a(n9006), .b(n7388) );
no02f01  g4206 ( .o(n9694), .a(n9693), .b(n9005) );
no02f01  g4207 ( .o(n2409), .a(n9694), .b(n9011) );
in01f01  g4208 ( .o(n9696), .a(net_10176) );
oa22f01  g4209 ( .o(n2419), .a(n7956), .b(n5597_1), .c(n7955), .d(n9696) );
no02f01  g4210 ( .o(n9698), .a(_net_10030), .b(n9024) );
no02f01  g4211 ( .o(n9699), .a(n7412), .b(_net_10460) );
in01f01  g4212 ( .o(n9700), .a(n9699) );
no02f01  g4213 ( .o(n9701), .a(n9025), .b(_net_10029) );
ao12f01  g4214 ( .o(n9702), .a(n9698), .b(n9701), .c(n9700) );
no02f01  g4215 ( .o(n9703), .a(_net_10459), .b(n5897) );
no02f01  g4216 ( .o(n9704), .a(_net_10027), .b(n9018) );
no02f01  g4217 ( .o(n9705), .a(_net_10028), .b(n9017) );
no02f01  g4218 ( .o(n9706), .a(n9705), .b(n9704) );
no02f01  g4219 ( .o(n9707), .a(n7389_1), .b(_net_10457) );
na02f01  g4220 ( .o(n9708), .a(n7396), .b(_net_10456) );
no02f01  g4221 ( .o(n9709), .a(_net_10455), .b(n7399) );
no02f01  g4222 ( .o(n9710), .a(n7396), .b(_net_10456) );
oa12f01  g4223 ( .o(n9711), .a(n9708), .b(n9710), .c(n9709) );
in01f01  g4224 ( .o(n9712), .a(n9711) );
no02f01  g4225 ( .o(n9713), .a(n9712), .b(n9707) );
in01f01  g4226 ( .o(n9714), .a(n9713) );
ao22f01  g4227 ( .o(n9715), .a(n9714), .b(n9706), .c(_net_10028), .d(n9017) );
in01f01  g4228 ( .o(n9716), .a(n9715) );
no02f01  g4229 ( .o(n9717), .a(n9716), .b(n9703) );
na02f01  g4230 ( .o(n9718), .a(n9717), .b(n9700) );
no02f01  g4231 ( .o(n9719), .a(n7379_1), .b(_net_10461) );
no02f01  g4232 ( .o(n9720), .a(_net_10031), .b(n9036) );
no02f01  g4233 ( .o(n9721), .a(n9720), .b(n9719) );
in01f01  g4234 ( .o(n9722), .a(n9721) );
ao12f01  g4235 ( .o(n9723), .a(n9722), .b(n9718), .c(n9702) );
na03f01  g4236 ( .o(n9724), .a(n9722), .b(n9718), .c(n9702) );
na02f01  g4237 ( .o(n9725), .a(n9724), .b(n7431) );
no02f01  g4238 ( .o(n9726), .a(n9014), .b(n9013) );
in01f01  g4239 ( .o(n9727), .a(n9726) );
no02f01  g4240 ( .o(n9728), .a(n9727), .b(n9018) );
in01f01  g4241 ( .o(n9729), .a(n9728) );
no02f01  g4242 ( .o(n9730), .a(n9729), .b(n9017) );
in01f01  g4243 ( .o(n9731), .a(n9730) );
no02f01  g4244 ( .o(n9732), .a(n9731), .b(n9033) );
na02f01  g4245 ( .o(n9733), .a(n9732), .b(_net_10461) );
no02f01  g4246 ( .o(n9734), .a(n9732), .b(_net_10461) );
no02f01  g4247 ( .o(n9735), .a(n9734), .b(n7451_1) );
ao22f01  g4248 ( .o(n9736), .a(n9735), .b(n9733), .c(n7453), .d(_net_10461) );
oa12f01  g4249 ( .o(n2424), .a(n9736), .b(n9725), .c(n9723) );
na04f01  g4250 ( .o(n9738), .a(n8021_1), .b(_net_9178), .c(net_9184), .d(_net_9183) );
no04f01  g4251 ( .o(n2429), .a(n9738), .b(n8027), .c(n8028), .d(_net_9177) );
in01f01  g4252 ( .o(n3146), .a(_net_10114) );
na02f01  g4253 ( .o(n9741), .a(n3146), .b(_net_10115) );
na02f01  g4254 ( .o(n9742), .a(_net_10114), .b(n7780) );
na02f01  g4255 ( .o(n2434), .a(n9742), .b(n9741) );
oa22f01  g4256 ( .o(n2444), .a(n7480_1), .b(n6773_1), .c(n7478), .d(n5585_1) );
in01f01  g4257 ( .o(n9745), .a(net_9585) );
no02f01  g4258 ( .o(n2458), .a(_net_9606), .b(n9745) );
in01f01  g4259 ( .o(n9747), .a(net_10506) );
na02f01  g4260 ( .o(n9748), .a(net_10490), .b(net_264) );
ao12f01  g4261 ( .o(n2463), .a(n9667), .b(n9748), .c(n9747) );
in01f01  g4262 ( .o(n9750), .a(_net_9190) );
oa22f01  g4263 ( .o(n2468), .a(n8349_1), .b(n8025), .c(n8347), .d(n9750) );
na02f01  g4264 ( .o(n9752), .a(n6699_1), .b(n6689_1) );
na02f01  g4265 ( .o(n9753), .a(n9752), .b(n6701) );
oa22f01  g4266 ( .o(n2477), .a(n9753), .b(n6688), .c(n6685), .d(n6689_1) );
na02f01  g4267 ( .o(n9755), .a(n7907), .b(_net_9161) );
oa12f01  g4268 ( .o(n9756), .a(n8754), .b(n9755), .c(n7920) );
no02f01  g4269 ( .o(n9757), .a(n9756), .b(_net_9354) );
in01f01  g4270 ( .o(n9758), .a(n9756) );
in01f01  g4271 ( .o(n9759), .a(n7921_1) );
na02f01  g4272 ( .o(n9760), .a(n7896), .b(x6599) );
no03f01  g4273 ( .o(n9761), .a(n9760), .b(n9759), .c(n7908) );
no02f01  g4274 ( .o(n9762), .a(n7889_1), .b(n7732) );
oa12f01  g4275 ( .o(n9763), .a(n9761), .b(n9762), .c(n9758) );
na03f01  g4276 ( .o(n9764), .a(n7895), .b(_net_9354), .c(n7888) );
na02f01  g4277 ( .o(n9765), .a(_net_9356), .b(x6599) );
oa22f01  g4278 ( .o(n9766), .a(n9765), .b(n8754), .c(n9764), .d(n5658) );
in01f01  g4279 ( .o(n9767), .a(_net_9355) );
no02f01  g4280 ( .o(n9768), .a(n9767), .b(n5658) );
na02f01  g4281 ( .o(n9769), .a(n9768), .b(n7887) );
oa12f01  g4282 ( .o(n9770), .a(_net_9354), .b(n8754), .c(net_9151) );
in01f01  g4283 ( .o(n9771), .a(_net_9353) );
no02f01  g4284 ( .o(n9772), .a(n9771), .b(n5658) );
na02f01  g4285 ( .o(n9773), .a(n7885_1), .b(n7889_1) );
no03f01  g4286 ( .o(n9774), .a(n9765), .b(n7732), .c(_net_9160) );
ao22f01  g4287 ( .o(n9775), .a(n9774), .b(_net_9354), .c(n9773), .d(n9772) );
oa12f01  g4288 ( .o(n9776), .a(n9775), .b(n9770), .c(n9769) );
ao12f01  g4289 ( .o(n9777), .a(n9776), .b(n9766), .c(n9762) );
oa12f01  g4290 ( .o(n2482), .a(n9777), .b(n9763), .c(n9757) );
no02f01  g4291 ( .o(n9779), .a(n7032), .b(n7028) );
na02f01  g4292 ( .o(n9780), .a(n9779), .b(n7030_1) );
in01f01  g4293 ( .o(n9781), .a(n7030_1) );
oa12f01  g4294 ( .o(n9782), .a(n9781), .b(n7032), .c(n7028) );
na02f01  g4295 ( .o(n2487), .a(n9782), .b(n9780) );
in01f01  g4296 ( .o(n9784), .a(net_9947) );
oa22f01  g4297 ( .o(n2492), .a(n5694), .b(n9784), .c(n5692), .d(n5597_1) );
in01f01  g4298 ( .o(n9786), .a(_net_9642) );
no03f01  g4299 ( .o(n9787), .a(n9540), .b(n7966), .c(n9786) );
no02f01  g4300 ( .o(n9788), .a(n9550), .b(n8756) );
no02f01  g4301 ( .o(n9789), .a(n8752), .b(n9786) );
oa12f01  g4302 ( .o(n9790), .a(_net_9641), .b(n9789), .c(n9788) );
in01f01  g4303 ( .o(n9791), .a(n9496) );
na02f01  g4304 ( .o(n9792), .a(n9545), .b(_net_9642) );
oa22f01  g4305 ( .o(n9793), .a(n9792), .b(n8773), .c(n9791), .d(n9786) );
ao12f01  g4306 ( .o(n9794), .a(n9793), .b(n9495), .c(_net_9642) );
oa12f01  g4307 ( .o(n9795), .a(n9794), .b(n9790), .c(n9490) );
no02f01  g4308 ( .o(n9796), .a(n9795), .b(n9787) );
no02f01  g4309 ( .o(n2502), .a(n9796), .b(n9500) );
in01f01  g4310 ( .o(n9798), .a(net_10192) );
no04f01  g4311 ( .o(n9799), .a(n5935_1), .b(n8579), .c(n8578), .d(_net_9563) );
na02f01  g4312 ( .o(n9800), .a(n9799), .b(net_10175) );
ao12f01  g4313 ( .o(n2507), .a(n8577_1), .b(n9800), .c(n9798) );
no02f01  g4314 ( .o(n9802), .a(n5918), .b(_net_187) );
no02f01  g4315 ( .o(n9803), .a(_net_9609), .b(_net_9608) );
in01f01  g4316 ( .o(n9804), .a(net_9610) );
na03f01  g4317 ( .o(n9805), .a(n9803), .b(n5921_1), .c(n9804) );
ao12f01  g4318 ( .o(n9806), .a(net_9607), .b(n9805), .c(n7725) );
ao12f01  g4319 ( .o(n9807), .a(n9806), .b(n9803), .c(n9802) );
no03f01  g4320 ( .o(n2512), .a(n9807), .b(n6460_1), .c(n7970) );
no02f01  g4321 ( .o(n2517), .a(n6164_1), .b(n6174) );
no02f01  g4322 ( .o(n9810), .a(n8814_1), .b(n7073_1) );
in01f01  g4323 ( .o(n9811), .a(n9810) );
no02f01  g4324 ( .o(n9812), .a(n9811), .b(n7605_1) );
in01f01  g4325 ( .o(n9813), .a(n9812) );
no02f01  g4326 ( .o(n9814), .a(n9813), .b(n8469) );
in01f01  g4327 ( .o(n9815), .a(n9814) );
no02f01  g4328 ( .o(n9816), .a(n9815), .b(n7545) );
in01f01  g4329 ( .o(n9817), .a(n9816) );
no02f01  g4330 ( .o(n9818), .a(n9817), .b(n7552_1) );
in01f01  g4331 ( .o(n9819), .a(n9818) );
no02f01  g4332 ( .o(n9820), .a(n9819), .b(n7536) );
na02f01  g4333 ( .o(n9821), .a(n9820), .b(_net_9299) );
ao12f01  g4334 ( .o(n9822), .a(n8810), .b(n9821), .c(n7516) );
oa12f01  g4335 ( .o(n9823), .a(n9822), .b(n9821), .c(n7516) );
oa12f01  g4336 ( .o(n2522), .a(n9823), .b(n8817), .c(n7516) );
in01f01  g4337 ( .o(n9825), .a(net_9846) );
in01f01  g4338 ( .o(n9826), .a(net_9838) );
no02f01  g4339 ( .o(n9827), .a(n6973), .b(n9826) );
no02f01  g4340 ( .o(n9828), .a(n9827), .b(n7477) );
no02f01  g4341 ( .o(n9829), .a(n9828), .b(n5658) );
oa12f01  g4342 ( .o(n9830), .a(n9829), .b(n7479), .c(x4587) );
na02f01  g4343 ( .o(n9831), .a(n9828), .b(x6599) );
oa12f01  g4344 ( .o(n2527), .a(n9830), .b(n9831), .c(n9825) );
na02f01  g4345 ( .o(n9833), .a(n8202), .b(_net_10351) );
na02f01  g4346 ( .o(n9834), .a(n9129), .b(n9128) );
na03f01  g4347 ( .o(n9835), .a(n9834), .b(n9131), .c(n8200_1) );
in01f01  g4348 ( .o(n9836), .a(n9095) );
in01f01  g4349 ( .o(n9837), .a(n9096) );
na03f01  g4350 ( .o(n9838), .a(n9837), .b(n9836), .c(n9094) );
in01f01  g4351 ( .o(n9839), .a(n9094) );
oa12f01  g4352 ( .o(n9840), .a(n9095), .b(n9096), .c(n9839) );
na03f01  g4353 ( .o(n9841), .a(n9840), .b(n9838), .c(n8183) );
na03f01  g4354 ( .o(n2541), .a(n9841), .b(n9835), .c(n9833) );
in01f01  g4355 ( .o(n9843), .a(net_9584) );
na02f01  g4356 ( .o(n9844), .a(_net_177), .b(n9843) );
oa22f01  g4357 ( .o(n9845), .a(n7573), .b(net_9576), .c(n7071), .d(net_9577) );
in01f01  g4358 ( .o(n9846), .a(net_9575) );
in01f01  g4359 ( .o(n9847), .a(net_9574) );
ao12f01  g4360 ( .o(n9848), .a(n9846), .b(n9847), .c(_net_167) );
na03f01  g4361 ( .o(n9849), .a(n9847), .b(_net_167), .c(n9846) );
ao12f01  g4362 ( .o(n9850), .a(n9848), .b(n9849), .c(n5916) );
no02f01  g4363 ( .o(n9851), .a(n9850), .b(n9845) );
in01f01  g4364 ( .o(n9852), .a(net_9576) );
no03f01  g4365 ( .o(n9853), .a(_net_169), .b(_net_170), .c(n9852) );
in01f01  g4366 ( .o(n9854), .a(net_9577) );
na02f01  g4367 ( .o(n9855), .a(n7573), .b(net_9577) );
oa22f01  g4368 ( .o(n9856), .a(n9855), .b(n9852), .c(_net_170), .d(n9854) );
no03f01  g4369 ( .o(n9857), .a(n9856), .b(n9853), .c(n9851) );
oa22f01  g4370 ( .o(n9858), .a(n8466), .b(_net_9580), .c(n7554), .d(_net_9581) );
oa22f01  g4371 ( .o(n9859), .a(n8468), .b(net_9578), .c(n5975), .d(net_9579) );
no03f01  g4372 ( .o(n9860), .a(n9859), .b(n9858), .c(n9857) );
in01f01  g4373 ( .o(n9861), .a(net_9578) );
no03f01  g4374 ( .o(n9862), .a(_net_171), .b(_net_172), .c(n9861) );
in01f01  g4375 ( .o(n9863), .a(net_9579) );
no03f01  g4376 ( .o(n9864), .a(_net_171), .b(n9863), .c(n9861) );
no02f01  g4377 ( .o(n9865), .a(_net_172), .b(n9863) );
no03f01  g4378 ( .o(n9866), .a(n9865), .b(n9864), .c(n9862) );
no02f01  g4379 ( .o(n9867), .a(n9866), .b(n9858) );
in01f01  g4380 ( .o(n9868), .a(_net_9581) );
in01f01  g4381 ( .o(n9869), .a(_net_9580) );
no03f01  g4382 ( .o(n9870), .a(_net_173), .b(n9869), .c(n9868) );
na02f01  g4383 ( .o(n9871), .a(n7554), .b(_net_9580) );
oa22f01  g4384 ( .o(n9872), .a(n9871), .b(_net_173), .c(_net_174), .d(n9868) );
no04f01  g4385 ( .o(n9873), .a(n9872), .b(n9870), .c(n9867), .d(n9860) );
oa22f01  g4386 ( .o(n9874), .a(n5990), .b(net_9583), .c(n5989), .d(net_9582) );
in01f01  g4387 ( .o(n9875), .a(net_9583) );
in01f01  g4388 ( .o(n9876), .a(net_9582) );
no03f01  g4389 ( .o(n9877), .a(_net_175), .b(n9876), .c(n9875) );
no03f01  g4390 ( .o(n9878), .a(_net_176), .b(_net_175), .c(n9876) );
oa22f01  g4391 ( .o(n9879), .a(_net_177), .b(n9843), .c(_net_176), .d(n9875) );
no03f01  g4392 ( .o(n9880), .a(n9879), .b(n9878), .c(n9877) );
oa12f01  g4393 ( .o(n9881), .a(n9880), .b(n9874), .c(n9873) );
in01f01  g4394 ( .o(n9882), .a(net_9587) );
no02f01  g4395 ( .o(n9883), .a(net_9586), .b(net_9585) );
na02f01  g4396 ( .o(n9884), .a(n9883), .b(n9882) );
ao12f01  g4397 ( .o(n2546), .a(n9884), .b(n9881), .c(n9844) );
oa22f01  g4398 ( .o(n2551), .a(n5694), .b(n5706), .c(n5692), .d(n5540) );
ao22f01  g4399 ( .o(n9887), .a(n5842), .b(net_9700), .c(n5841), .d(net_140) );
na02f01  g4400 ( .o(n9888), .a(n5847), .b(net_9997) );
ao22f01  g4401 ( .o(n9889), .a(n5850), .b(net_9799), .c(n5849_1), .d(net_9898) );
na03f01  g4402 ( .o(n2556), .a(n9889), .b(n9888), .c(n9887) );
no02f01  g4403 ( .o(n9891), .a(n8703), .b(net_9652) );
no03f01  g4404 ( .o(n2564), .a(n9891), .b(n9603), .c(net_9151) );
no02f01  g4405 ( .o(n9893), .a(n9074), .b(_net_10228) );
in01f01  g4406 ( .o(n9894), .a(n9893) );
na02f01  g4407 ( .o(n9895), .a(n9074), .b(_net_10228) );
na02f01  g4408 ( .o(n2572), .a(n9895), .b(n9894) );
ao12f01  g4409 ( .o(n9897), .a(n5658), .b(n6532), .c(net_248) );
ao22f01  g4410 ( .o(n9898), .a(n6535), .b(x5003), .c(n6534), .d(net_10008) );
na02f01  g4411 ( .o(n2577), .a(n9898), .b(n9897) );
in01f01  g4412 ( .o(n9900), .a(_net_10318) );
ao12f01  g4413 ( .o(n9901), .a(n5658), .b(n5774), .c(x5289) );
oa12f01  g4414 ( .o(n2582), .a(n9901), .b(n5770), .c(n9900) );
no02f01  g4415 ( .o(n9903), .a(n6686), .b(net_9227) );
in01f01  g4416 ( .o(n9904), .a(n9903) );
in01f01  g4417 ( .o(n9905), .a(net_9223) );
in01f01  g4418 ( .o(n9906), .a(net_9222) );
in01f01  g4419 ( .o(n9907), .a(net_9221) );
in01f01  g4420 ( .o(n9908), .a(net_9220) );
in01f01  g4421 ( .o(n9909), .a(net_9219) );
no02f01  g4422 ( .o(n9910), .a(n9909), .b(n9908) );
in01f01  g4423 ( .o(n9911), .a(n9910) );
no02f01  g4424 ( .o(n9912), .a(n9911), .b(n9907) );
in01f01  g4425 ( .o(n9913), .a(n9912) );
no02f01  g4426 ( .o(n9914), .a(n9913), .b(n9906) );
in01f01  g4427 ( .o(n9915), .a(n9914) );
no02f01  g4428 ( .o(n9916), .a(n9915), .b(n9905) );
no02f01  g4429 ( .o(n9917), .a(n9916), .b(net_9224) );
in01f01  g4430 ( .o(n9918), .a(net_9224) );
in01f01  g4431 ( .o(n9919), .a(n9916) );
no02f01  g4432 ( .o(n9920), .a(n9919), .b(n9918) );
no03f01  g4433 ( .o(n2587), .a(n9920), .b(n9917), .c(n9904) );
na02f01  g4434 ( .o(n9922), .a(n7937), .b(net_258) );
na02f01  g4435 ( .o(n9923), .a(n7936), .b(net_9788) );
ao22f01  g4436 ( .o(n9924), .a(n7943), .b(_net_10227), .c(n7942), .d(x4209) );
na04f01  g4437 ( .o(n2592), .a(n9924), .b(n9923), .c(n9922), .d(n7939) );
na02f01  g4438 ( .o(n9926), .a(n8202), .b(_net_10363) );
no02f01  g4439 ( .o(n9927), .a(n7029), .b(n7031) );
oa12f01  g4440 ( .o(n9928), .a(n8200_1), .b(n9927), .c(n8187) );
in01f01  g4441 ( .o(n9929), .a(n8168) );
na03f01  g4442 ( .o(n9930), .a(n8171), .b(n8169), .c(n9929) );
in01f01  g4443 ( .o(n9931), .a(n8169) );
oa12f01  g4444 ( .o(n9932), .a(n9931), .b(n8170_1), .c(n8168) );
na03f01  g4445 ( .o(n9933), .a(n9932), .b(n9930), .c(n8183) );
na03f01  g4446 ( .o(n2597), .a(n9933), .b(n9928), .c(n9926) );
na02f01  g4447 ( .o(n9935), .a(n6056), .b(_net_232) );
na02f01  g4448 ( .o(n9936), .a(n6055), .b(net_9960) );
ao22f01  g4449 ( .o(n9937), .a(n6062_1), .b(x6028), .c(n6060), .d(_net_10411) );
na04f01  g4450 ( .o(n2602), .a(n9937), .b(n9936), .c(n9935), .d(n6058) );
in01f01  g4451 ( .o(n9939), .a(x3733) );
in01f01  g4452 ( .o(n9940), .a(_net_10348) );
na02f01  g4453 ( .o(n9941), .a(_net_10349), .b(n9940) );
ao12f01  g4454 ( .o(n2607), .a(n5658), .b(n9941), .c(n9939) );
in01f01  g4455 ( .o(n9943), .a(_net_9950) );
no02f01  g4456 ( .o(n9944), .a(n9943), .b(_net_9949) );
in01f01  g4457 ( .o(n9945), .a(n9944) );
no03f01  g4458 ( .o(n9946), .a(_net_10365), .b(_net_10370), .c(_net_10372) );
na03f01  g4459 ( .o(n9947), .a(n9946), .b(n6996), .c(n9321) );
no04f01  g4460 ( .o(n9948), .a(_net_10367), .b(_net_10369), .c(_net_10366), .d(_net_10368) );
na02f01  g4461 ( .o(n9949), .a(n9948), .b(n7024) );
no02f01  g4462 ( .o(n9950), .a(n9949), .b(n9947) );
no02f01  g4463 ( .o(n2612), .a(n9950), .b(n9945) );
ao22f01  g4464 ( .o(n9952), .a(n5842), .b(net_9725), .c(n5841), .d(_net_165) );
na02f01  g4465 ( .o(n9953), .a(n5847), .b(net_10022) );
ao22f01  g4466 ( .o(n9954), .a(n5850), .b(net_9824), .c(n5849_1), .d(net_9923) );
na03f01  g4467 ( .o(n2617), .a(n9954), .b(n9953), .c(n9952) );
in01f01  g4468 ( .o(n9956), .a(net_9544) );
oa12f01  g4469 ( .o(n2622), .a(n9956), .b(n5739_1), .c(n5738) );
na02f01  g4470 ( .o(n9958), .a(n8079), .b(_net_10529) );
no04f01  g4471 ( .o(n2627), .a(n9958), .b(n6559), .c(n5660), .d(x6496) );
na02f01  g4472 ( .o(n9960), .a(n6349), .b(n6245) );
oa22f01  g4473 ( .o(n2632), .a(n9960), .b(n6348), .c(n6349), .d(n8853_1) );
no02f01  g4474 ( .o(n2637), .a(n7703), .b(net_9228) );
ao22f01  g4475 ( .o(n9963), .a(n5842), .b(net_9748), .c(n5841), .d(_net_184) );
na02f01  g4476 ( .o(n9964), .a(n5847), .b(net_10045) );
ao22f01  g4477 ( .o(n9965), .a(n5850), .b(net_9847), .c(n5849_1), .d(net_9946) );
na03f01  g4478 ( .o(n2642), .a(n9965), .b(n9964), .c(n9963) );
in01f01  g4479 ( .o(n9967), .a(_net_10101) );
ao12f01  g4480 ( .o(n9968), .a(n5658), .b(n6160_1), .c(x5722) );
oa12f01  g4481 ( .o(n2652), .a(n9968), .b(n6159), .c(n9967) );
ao22f01  g4482 ( .o(n9970), .a(n5842), .b(net_9747), .c(n5841), .d(_net_183) );
na02f01  g4483 ( .o(n9971), .a(n5847), .b(net_10044) );
ao22f01  g4484 ( .o(n9972), .a(n5850), .b(net_9846), .c(n5849_1), .d(net_9945) );
na03f01  g4485 ( .o(n2657), .a(n9972), .b(n9971), .c(n9970) );
ao22f01  g4486 ( .o(n9974), .a(n6602), .b(net_10004), .c(n6597), .d(net_9739) );
ao22f01  g4487 ( .o(n9975), .a(n6577), .b(net_9675), .c(n6555), .d(net_9972) );
in01f01  g4488 ( .o(n9976), .a(net_9937) );
in01f01  g4489 ( .o(n9977), .a(net_9806) );
in01f01  g4490 ( .o(n9978), .a(n6580) );
oa22f01  g4491 ( .o(n9979), .a(n6966_1), .b(n9976), .c(n9978), .d(n9977) );
na02f01  g4492 ( .o(n9980), .a(n6585), .b(net_9707) );
na02f01  g4493 ( .o(n9981), .a(n6582), .b(net_9905) );
na02f01  g4494 ( .o(n9982), .a(n9981), .b(n9980) );
ao22f01  g4495 ( .o(n9983), .a(n6590), .b(net_10036), .c(n6573), .d(net_9873) );
ao22f01  g4496 ( .o(n9984), .a(n6599_1), .b(net_9838), .c(n6584_1), .d(net_9774) );
na02f01  g4497 ( .o(n9985), .a(n9984), .b(n9983) );
no03f01  g4498 ( .o(n9986), .a(n9985), .b(n9982), .c(n9979) );
na03f01  g4499 ( .o(n2667), .a(n9986), .b(n9975), .c(n9974) );
ao12f01  g4500 ( .o(n9988), .a(n5658), .b(n6875_1), .c(net_237) );
ao22f01  g4501 ( .o(n9989), .a(n6878), .b(x5722), .c(n6877), .d(net_9898) );
na02f01  g4502 ( .o(n2671), .a(n9989), .b(n9988) );
na02f01  g4503 ( .o(n9991), .a(n6349), .b(n6254_1) );
oa22f01  g4504 ( .o(n2676), .a(n9991), .b(n6348), .c(n6349), .d(n8860) );
in01f01  g4505 ( .o(n9993), .a(n7040) );
no03f01  g4506 ( .o(n9994), .a(n7050), .b(n7047), .c(n9993) );
in01f01  g4507 ( .o(n9995), .a(n9994) );
no02f01  g4508 ( .o(n9996), .a(n7051), .b(n7006) );
in01f01  g4509 ( .o(n9997), .a(n9996) );
na02f01  g4510 ( .o(n9998), .a(n9997), .b(n9995) );
na02f01  g4511 ( .o(n9999), .a(n9996), .b(n9994) );
na02f01  g4512 ( .o(n2681), .a(n9999), .b(n9998) );
in01f01  g4513 ( .o(n10001), .a(net_9275) );
na02f01  g4514 ( .o(n10002), .a(n10001), .b(net_9274) );
in01f01  g4515 ( .o(n10003), .a(net_9274) );
na02f01  g4516 ( .o(n10004), .a(net_9275), .b(n10003) );
na03f01  g4517 ( .o(n10005), .a(n5914), .b(n7754), .c(x6599) );
ao12f01  g4518 ( .o(n2695), .a(n10005), .b(n10004), .c(n10002) );
na02f01  g4519 ( .o(n10007), .a(n8202), .b(_net_10352) );
na02f01  g4520 ( .o(n10008), .a(n9131), .b(n9087) );
na03f01  g4521 ( .o(n10009), .a(n10008), .b(n9133), .c(n8200_1) );
no02f01  g4522 ( .o(n10010), .a(n9093), .b(n9088) );
in01f01  g4523 ( .o(n10011), .a(n10010) );
na02f01  g4524 ( .o(n10012), .a(n10011), .b(n9098) );
na02f01  g4525 ( .o(n10013), .a(n10010), .b(n9097) );
na03f01  g4526 ( .o(n10014), .a(n10013), .b(n10012), .c(n8183) );
na03f01  g4527 ( .o(n2700), .a(n10014), .b(n10009), .c(n10007) );
no02f01  g4528 ( .o(n10016), .a(net_9219), .b(net_9220) );
no03f01  g4529 ( .o(n2705), .a(n10016), .b(n9910), .c(n9904) );
ao22f01  g4530 ( .o(n10018), .a(n5842), .b(net_9705), .c(n5841), .d(net_145) );
na02f01  g4531 ( .o(n10019), .a(n5847), .b(net_10002) );
ao22f01  g4532 ( .o(n10020), .a(n5850), .b(net_9804), .c(n5849_1), .d(net_9903) );
na03f01  g4533 ( .o(n2710), .a(n10020), .b(n10019), .c(n10018) );
in01f01  g4534 ( .o(n10022), .a(net_10494) );
oa22f01  g4535 ( .o(n2715), .a(n7467), .b(n5637), .c(n7465_1), .d(n10022) );
ao12f01  g4536 ( .o(n10024), .a(n5658), .b(n6532), .c(net_251) );
ao22f01  g4537 ( .o(n10025), .a(n6535), .b(x4781), .c(n6534), .d(net_10011) );
na02f01  g4538 ( .o(n2725), .a(n10025), .b(n10024) );
na02f01  g4539 ( .o(n10027), .a(n6172), .b(_net_10219) );
na02f01  g4540 ( .o(n2730), .a(n10027), .b(n8963) );
ao22f01  g4541 ( .o(n10029), .a(n5842), .b(net_9679), .c(n5841), .d(_net_117) );
na02f01  g4542 ( .o(n10030), .a(n5847), .b(net_9976) );
ao22f01  g4543 ( .o(n10031), .a(n5850), .b(net_9778), .c(n5849_1), .d(net_9877) );
na03f01  g4544 ( .o(n2735), .a(n10031), .b(n10030), .c(n10029) );
ao22f01  g4545 ( .o(n10033), .a(n5842), .b(net_9755), .c(n5841), .d(_net_191) );
na02f01  g4546 ( .o(n10034), .a(n5847), .b(net_10052) );
ao22f01  g4547 ( .o(n10035), .a(n5850), .b(net_9854), .c(n5849_1), .d(net_9953) );
na03f01  g4548 ( .o(n2745), .a(n10035), .b(n10034), .c(n10033) );
ao22f01  g4549 ( .o(n10037), .a(n5743), .b(x1418), .c(n5742), .d(_net_9420) );
oa12f01  g4550 ( .o(n2750), .a(n10037), .b(n5741), .c(n9409) );
ao12f01  g4551 ( .o(n10039), .a(n5658), .b(n6052_1), .c(x4285) );
oa12f01  g4552 ( .o(n2755), .a(n10039), .b(n6048), .c(n9027) );
oa22f01  g4553 ( .o(n2760), .a(n5907), .b(n9055), .c(n5905), .d(n5609) );
in01f01  g4554 ( .o(n10042), .a(n8106_1) );
no02f01  g4555 ( .o(n10043), .a(n8105), .b(n5658) );
in01f01  g4556 ( .o(n10044), .a(n10043) );
no02f01  g4557 ( .o(n10045), .a(n10044), .b(n10042) );
oa12f01  g4558 ( .o(n10046), .a(n10045), .b(n7446), .c(_net_9383) );
ao12f01  g4559 ( .o(n10047), .a(n5658), .b(n6142), .c(n8104) );
na03f01  g4560 ( .o(n10048), .a(n10047), .b(n6136_1), .c(_net_9383) );
na03f01  g4561 ( .o(n10049), .a(n6140), .b(_net_9383), .c(x6599) );
na03f01  g4562 ( .o(n2765), .a(n10049), .b(n10048), .c(n10046) );
no02f01  g4563 ( .o(n10051), .a(n6687), .b(_net_9201) );
ao12f01  g4564 ( .o(n2774), .a(n10051), .b(n6685), .c(_net_9201) );
oa22f01  g4565 ( .o(n2779), .a(n7367), .b(n5786), .c(n7365_1), .d(n5640) );
oa22f01  g4566 ( .o(n2784), .a(n5907), .b(n7379_1), .c(n5905), .d(n5606) );
no03f01  g4567 ( .o(n10055), .a(n6474_1), .b(n6489_1), .c(n6463) );
no02f01  g4568 ( .o(n10056), .a(n6502), .b(n6489_1) );
na02f01  g4569 ( .o(n10057), .a(n10056), .b(_net_9248) );
no02f01  g4570 ( .o(n10058), .a(n6511), .b(n6489_1) );
ao22f01  g4571 ( .o(n10059), .a(n10058), .b(n6860), .c(n6500), .d(_net_9241) );
na02f01  g4572 ( .o(n10060), .a(n10059), .b(n10057) );
na03f01  g4573 ( .o(n10061), .a(n6850), .b(n6486), .c(_net_9241) );
in01f01  g4574 ( .o(n10062), .a(n6136) );
ao12f01  g4575 ( .o(n10063), .a(n6491), .b(n10062), .c(n6489_1) );
no02f01  g4576 ( .o(n10064), .a(n6477), .b(n6489_1) );
no03f01  g4577 ( .o(n10065), .a(_net_9209), .b(n6520), .c(n6489_1) );
no04f01  g4578 ( .o(n10066), .a(n10065), .b(n10064), .c(n10063), .d(n6490) );
oa12f01  g4579 ( .o(n10067), .a(n10056), .b(n6508), .c(n6506) );
na03f01  g4580 ( .o(n10068), .a(n10067), .b(n10066), .c(n10061) );
no03f01  g4581 ( .o(n10069), .a(n10068), .b(n10060), .c(n10055) );
no02f01  g4582 ( .o(n2789), .a(n10069), .b(n6526_1) );
ao22f01  g4583 ( .o(n10071), .a(n5842), .b(net_9668), .c(n5841), .d(net_106) );
na02f01  g4584 ( .o(n10072), .a(n5847), .b(net_9965) );
ao22f01  g4585 ( .o(n10073), .a(n5850), .b(net_9767), .c(n5849_1), .d(net_9866) );
na03f01  g4586 ( .o(n2803), .a(n10073), .b(n10072), .c(n10071) );
ao22f01  g4587 ( .o(n10075), .a(n5842), .b(net_9665), .c(n5841), .d(net_103) );
na02f01  g4588 ( .o(n10076), .a(n5847), .b(net_9962) );
ao22f01  g4589 ( .o(n10077), .a(n5850), .b(net_9764), .c(n5849_1), .d(net_9863) );
na03f01  g4590 ( .o(n2808), .a(n10077), .b(n10076), .c(n10075) );
na02f01  g4591 ( .o(n10079), .a(n6038), .b(net_252) );
na02f01  g4592 ( .o(n10080), .a(n6037_1), .b(net_9881) );
ao22f01  g4593 ( .o(n10081), .a(n6044), .b(x4694), .c(n6042_1), .d(_net_10326) );
na04f01  g4594 ( .o(n2813), .a(n10081), .b(n10080), .c(n10079), .d(n6040) );
in01f01  g4595 ( .o(n10083), .a(net_10507) );
na02f01  g4596 ( .o(n10084), .a(n9799), .b(net_10490) );
ao12f01  g4597 ( .o(n2822), .a(n9667), .b(n10084), .c(n10083) );
no02f01  g4598 ( .o(n10086), .a(_net_9209), .b(n6520) );
in01f01  g4599 ( .o(n10087), .a(n10086) );
no02f01  g4600 ( .o(n10088), .a(n6502), .b(n6507_1) );
na03f01  g4601 ( .o(n10089), .a(n10088), .b(n6467), .c(n6853) );
ao12f01  g4602 ( .o(n10090), .a(n6507_1), .b(n10089), .c(n10087) );
na03f01  g4603 ( .o(n10091), .a(n6860), .b(_net_9236), .c(_net_9246) );
ao22f01  g4604 ( .o(n10092), .a(n10088), .b(_net_9248), .c(n6500), .d(_net_9246) );
na03f01  g4605 ( .o(n10093), .a(n6850), .b(n6486), .c(_net_9246) );
no02f01  g4606 ( .o(n10094), .a(net_9170), .b(_net_9246) );
no02f01  g4607 ( .o(n10095), .a(n10094), .b(n6475) );
ao12f01  g4608 ( .o(n10096), .a(n10095), .b(n6494), .c(_net_9246) );
na04f01  g4609 ( .o(n10097), .a(n10096), .b(n10093), .c(n10092), .d(n10091) );
na02f01  g4610 ( .o(n10098), .a(_net_9246), .b(_net_9238) );
ao22f01  g4611 ( .o(n10099), .a(n10088), .b(n6853), .c(n7747), .d(n6471) );
oa22f01  g4612 ( .o(n10100), .a(n10099), .b(n6504), .c(n10098), .d(n6474_1) );
no03f01  g4613 ( .o(n10101), .a(n10100), .b(n10097), .c(n10090) );
no02f01  g4614 ( .o(n2836), .a(n10101), .b(n6526_1) );
ao12f01  g4615 ( .o(n10103), .a(n5658), .b(n7844), .c(net_240) );
ao22f01  g4616 ( .o(n10104), .a(n7847), .b(x5548), .c(n7846), .d(net_9802) );
na02f01  g4617 ( .o(n2841), .a(n10104), .b(n10103) );
in01f01  g4618 ( .o(n10106), .a(n6492) );
ao12f01  g4619 ( .o(n10107), .a(n6511), .b(n6861_1), .c(n10106) );
no03f01  g4620 ( .o(n10108), .a(n7482), .b(n6485), .c(n6511) );
na03f01  g4621 ( .o(n10109), .a(_net_9240), .b(n6677), .c(_net_9236) );
no02f01  g4622 ( .o(n10110), .a(n6477), .b(n6511) );
ao12f01  g4623 ( .o(n10111), .a(n6489_1), .b(n6511), .c(n6480) );
no03f01  g4624 ( .o(n10112), .a(n6497), .b(_net_9169), .c(n6511) );
ao12f01  g4625 ( .o(n10113), .a(n6520), .b(n6864), .c(n6511) );
no04f01  g4626 ( .o(n10114), .a(n10113), .b(n10112), .c(n10111), .d(n10110) );
na03f01  g4627 ( .o(n10115), .a(n10114), .b(n10109), .c(n6851_1) );
no03f01  g4628 ( .o(n10116), .a(n10115), .b(n10108), .c(n10107) );
no03f01  g4629 ( .o(n10117), .a(n6474_1), .b(n6511), .c(n6463) );
na02f01  g4630 ( .o(n10118), .a(n6853), .b(_net_9236) );
no04f01  g4631 ( .o(n10119), .a(n10118), .b(n6505), .c(n6502), .d(n6504) );
ao12f01  g4632 ( .o(n10120), .a(n7852), .b(n6471), .c(n6511) );
no04f01  g4633 ( .o(n10121), .a(n10118), .b(n6502), .c(n6468), .d(n6507_1) );
no04f01  g4634 ( .o(n10122), .a(n10121), .b(n10120), .c(n10119), .d(n10117) );
ao12f01  g4635 ( .o(n2846), .a(n6526_1), .b(n10122), .c(n10116) );
in01f01  g4636 ( .o(n10124), .a(net_10072) );
oa22f01  g4637 ( .o(n2855), .a(n6989_1), .b(n5570), .c(n6988), .d(n10124) );
no02f01  g4638 ( .o(n10126), .a(_net_9246), .b(_net_9245) );
no02f01  g4639 ( .o(n10127), .a(_net_9244), .b(_net_9243) );
na04f01  g4640 ( .o(n10128), .a(n10127), .b(n10126), .c(n8446), .d(n6489_1) );
no02f01  g4641 ( .o(n10129), .a(n8451), .b(_net_9235) );
no02f01  g4642 ( .o(n10130), .a(_net_9236), .b(_net_9247) );
in01f01  g4643 ( .o(n10131), .a(n8452_1) );
ao12f01  g4644 ( .o(n10132), .a(n10131), .b(n7852), .c(n6851_1) );
na04f01  g4645 ( .o(n10133), .a(n10132), .b(n10130), .c(n10129), .d(n6863) );
oa12f01  g4646 ( .o(n10134), .a(n6491), .b(n10133), .c(n10128) );
na03f01  g4647 ( .o(n10135), .a(n6679_1), .b(n8509), .c(x494) );
ao12f01  g4648 ( .o(n2860), .a(n10135), .b(n10134), .c(n10106) );
in01f01  g4649 ( .o(n10137), .a(net_10295) );
na02f01  g4650 ( .o(n10138), .a(n8768), .b(net_10280) );
ao12f01  g4651 ( .o(n2864), .a(n5911), .b(n10138), .c(n10137) );
in01f01  g4652 ( .o(n10140), .a(_net_10361) );
no03f01  g4653 ( .o(n10141), .a(n9122), .b(_net_10360), .c(n10140) );
no02f01  g4654 ( .o(n10142), .a(n9122), .b(_net_10360) );
oa12f01  g4655 ( .o(n10143), .a(n8183), .b(n10142), .c(_net_10361) );
na02f01  g4656 ( .o(n10144), .a(n9142), .b(_net_10360) );
in01f01  g4657 ( .o(n10145), .a(n10144) );
na02f01  g4658 ( .o(n10146), .a(n10145), .b(_net_10361) );
ao12f01  g4659 ( .o(n10147), .a(n9144), .b(n10144), .c(n10140) );
ao22f01  g4660 ( .o(n10148), .a(n10147), .b(n10146), .c(n8202), .d(_net_10361) );
oa12f01  g4661 ( .o(n2869), .a(n10148), .b(n10143), .c(n10141) );
in01f01  g4662 ( .o(n10150), .a(x747) );
in01f01  g4663 ( .o(n10151), .a(net_9163) );
no02f01  g4664 ( .o(n10152), .a(n7446), .b(net_9289) );
no02f01  g4665 ( .o(n10153), .a(n10152), .b(net_8827) );
no02f01  g4666 ( .o(n10154), .a(n10153), .b(x3653) );
na02f01  g4667 ( .o(n10155), .a(n10154), .b(n10151) );
in01f01  g4668 ( .o(n10156), .a(n10154) );
na02f01  g4669 ( .o(n10157), .a(n10155), .b(n10156) );
no02f01  g4670 ( .o(n10158), .a(net_9289), .b(_net_9380) );
in01f01  g4671 ( .o(n10159), .a(n10158) );
no02f01  g4672 ( .o(n10160), .a(_net_9382), .b(_net_9383) );
no03f01  g4673 ( .o(n10161), .a(n10160), .b(n8107), .c(n6141_1) );
in01f01  g4674 ( .o(n10162), .a(n10161) );
no02f01  g4675 ( .o(n10163), .a(n10162), .b(n10159) );
in01f01  g4676 ( .o(n10164), .a(n6146) );
no02f01  g4677 ( .o(n10165), .a(n6763_1), .b(_net_9385) );
na02f01  g4678 ( .o(n10166), .a(n10165), .b(n6146) );
no02f01  g4679 ( .o(n10167), .a(n10161), .b(n10159) );
na02f01  g4680 ( .o(n10168), .a(n10167), .b(n10166) );
no02f01  g4681 ( .o(n10169), .a(n10168), .b(n10164) );
in01f01  g4682 ( .o(n10170), .a(n10169) );
no02f01  g4683 ( .o(n10171), .a(n10168), .b(n6146) );
in01f01  g4684 ( .o(n10172), .a(net_9269) );
in01f01  g4685 ( .o(n10173), .a(n10166) );
na02f01  g4686 ( .o(n10174), .a(n10167), .b(n10173) );
in01f01  g4687 ( .o(n10175), .a(_net_9309) );
no02f01  g4688 ( .o(n10176), .a(n10175), .b(net_9308) );
in01f01  g4689 ( .o(n10177), .a(net_9308) );
no02f01  g4690 ( .o(n10178), .a(_net_9309), .b(n10177) );
no02f01  g4691 ( .o(n10179), .a(n10178), .b(n10176) );
oa22f01  g4692 ( .o(n10180), .a(n10179), .b(n10158), .c(n10174), .d(n10172) );
ao12f01  g4693 ( .o(n10181), .a(n10180), .b(n10171), .c(n7104_1) );
oa12f01  g4694 ( .o(n10182), .a(n10181), .b(n10170), .c(net_9366) );
ao12f01  g4695 ( .o(n10183), .a(n10182), .b(n10163), .c(n7263) );
oa22f01  g4696 ( .o(n2874), .a(n10183), .b(n10157), .c(n10155), .d(n10150) );
ao22f01  g4697 ( .o(n10185), .a(n5842), .b(net_9741), .c(n5841), .d(_net_181) );
na02f01  g4698 ( .o(n10186), .a(n5847), .b(net_10038) );
ao22f01  g4699 ( .o(n10187), .a(n5850), .b(net_9840), .c(n5849_1), .d(net_9939) );
na03f01  g4700 ( .o(n2878), .a(n10187), .b(n10186), .c(n10185) );
oa22f01  g4701 ( .o(n2883), .a(n7367), .b(n5778), .c(n7365_1), .d(n5546) );
ao12f01  g4702 ( .o(n10190), .a(n5658), .b(n6875_1), .c(net_244) );
ao22f01  g4703 ( .o(n10191), .a(n6878), .b(x5289), .c(n6877), .d(net_9905) );
na02f01  g4704 ( .o(n2888), .a(n10191), .b(n10190) );
no02f01  g4705 ( .o(n10193), .a(n6774), .b(n6772) );
ao12f01  g4706 ( .o(n10194), .a(n6933), .b(n10193), .c(n6821_1) );
oa12f01  g4707 ( .o(n10195), .a(n10194), .b(n10193), .c(n6821_1) );
in01f01  g4708 ( .o(n10196), .a(n6841_1) );
no02f01  g4709 ( .o(n10197), .a(n6840), .b(_net_10253) );
no03f01  g4710 ( .o(n10198), .a(n10197), .b(n10196), .c(n6846_1) );
ao12f01  g4711 ( .o(n10199), .a(n10198), .b(n6168), .c(_net_10253) );
na02f01  g4712 ( .o(n2893), .a(n10199), .b(n10195) );
na02f01  g4713 ( .o(n10201), .a(n7672), .b(_net_10436) );
na02f01  g4714 ( .o(n2898), .a(n10201), .b(n7674) );
oa12f01  g4715 ( .o(n10203), .a(n6629_1), .b(n9150), .c(n6627) );
no02f01  g4716 ( .o(n10204), .a(n9150), .b(n6627) );
na02f01  g4717 ( .o(n10205), .a(n10204), .b(n9151) );
na02f01  g4718 ( .o(n2903), .a(n10205), .b(n10203) );
ao22f01  g4719 ( .o(n10207), .a(n5702), .b(x2333), .c(n5701), .d(_net_9404) );
oa12f01  g4720 ( .o(n2912), .a(n10207), .b(n5700_1), .c(n9409) );
in01f01  g4721 ( .o(n10209), .a(net_10393) );
no02f01  g4722 ( .o(n10210), .a(n7464), .b(n5769) );
na02f01  g4723 ( .o(n10211), .a(n7466), .b(n5689) );
oa22f01  g4724 ( .o(n2917), .a(n10211), .b(n5591), .c(n10210), .d(n10209) );
ao12f01  g4725 ( .o(n10213), .a(n5658), .b(n6875_1), .c(net_247) );
ao22f01  g4726 ( .o(n10214), .a(n6878), .b(x5077), .c(n6877), .d(net_9908) );
na02f01  g4727 ( .o(n2922), .a(n10214), .b(n10213) );
na02f01  g4728 ( .o(n10216), .a(n8032), .b(net_9181) );
na02f01  g4729 ( .o(n10217), .a(n8031_1), .b(n8025) );
na02f01  g4730 ( .o(n2927), .a(n10217), .b(n10216) );
ao12f01  g4731 ( .o(n10219), .a(n5658), .b(n6532), .c(net_242) );
ao22f01  g4732 ( .o(n10220), .a(n6535), .b(x5427), .c(n6534), .d(net_10002) );
na02f01  g4733 ( .o(n2932), .a(n10220), .b(n10219) );
oa22f01  g4734 ( .o(n2937), .a(n5907), .b(n7372), .c(n5905), .d(n5585_1) );
no02f01  g4735 ( .o(n10223), .a(n7059), .b(n7000) );
no02f01  g4736 ( .o(n10224), .a(n6997), .b(n6995) );
na02f01  g4737 ( .o(n10225), .a(n10224), .b(n10223) );
in01f01  g4738 ( .o(n10226), .a(n10224) );
oa12f01  g4739 ( .o(n10227), .a(n10226), .b(n7059), .c(n7000) );
na02f01  g4740 ( .o(n2946), .a(n10227), .b(n10225) );
oa12f01  g4741 ( .o(n10229), .a(n6641), .b(n6637), .c(n9524) );
in01f01  g4742 ( .o(n10230), .a(n10229) );
no02f01  g4743 ( .o(n10231), .a(n6643), .b(n6635) );
na02f01  g4744 ( .o(n10232), .a(n10231), .b(n10230) );
in01f01  g4745 ( .o(n10233), .a(n10231) );
na02f01  g4746 ( .o(n10234), .a(n10233), .b(n10229) );
na02f01  g4747 ( .o(n2951), .a(n10234), .b(n10232) );
oa22f01  g4748 ( .o(n2960), .a(n7480_1), .b(n6178), .c(n7478), .d(n5540) );
no02f01  g4749 ( .o(n10237), .a(_net_9370), .b(n7095_1) );
no02f01  g4750 ( .o(n10238), .a(n7110), .b(_net_9371) );
no02f01  g4751 ( .o(n10239), .a(n10238), .b(n10237) );
no02f01  g4752 ( .o(n10240), .a(n10239), .b(net_9369) );
na02f01  g4753 ( .o(n10241), .a(n10239), .b(net_9369) );
in01f01  g4754 ( .o(n10242), .a(n10241) );
no02f01  g4755 ( .o(n10243), .a(n7106), .b(_net_9372) );
no02f01  g4756 ( .o(n10244), .a(_net_9373), .b(n7097) );
no02f01  g4757 ( .o(n10245), .a(n10244), .b(n10243) );
no03f01  g4758 ( .o(n10246), .a(n10245), .b(n10242), .c(n10240) );
in01f01  g4759 ( .o(n10247), .a(n10240) );
in01f01  g4760 ( .o(n10248), .a(n10245) );
ao12f01  g4761 ( .o(n10249), .a(n10248), .b(n10241), .c(n10247) );
no02f01  g4762 ( .o(n10250), .a(_net_9374), .b(n7088) );
no02f01  g4763 ( .o(n10251), .a(n7104_1), .b(_net_9375) );
no02f01  g4764 ( .o(n10252), .a(n10251), .b(n10250) );
no02f01  g4765 ( .o(n10253), .a(_net_9376), .b(n6106) );
no02f01  g4766 ( .o(n10254), .a(n7089), .b(_net_9377) );
no03f01  g4767 ( .o(n10255), .a(n10254), .b(n10253), .c(n10252) );
in01f01  g4768 ( .o(n10256), .a(n10252) );
no02f01  g4769 ( .o(n10257), .a(n10254), .b(n10253) );
no02f01  g4770 ( .o(n10258), .a(n10257), .b(n10256) );
no02f01  g4771 ( .o(n10259), .a(n10258), .b(n10255) );
in01f01  g4772 ( .o(n10260), .a(n10259) );
no03f01  g4773 ( .o(n10261), .a(n10260), .b(n10249), .c(n10246) );
no02f01  g4774 ( .o(n10262), .a(n10249), .b(n10246) );
no02f01  g4775 ( .o(n10263), .a(n10259), .b(n10262) );
no02f01  g4776 ( .o(n10264), .a(n10263), .b(n10261) );
no02f01  g4777 ( .o(n10265), .a(n10264), .b(n7335) );
in01f01  g4778 ( .o(n10266), .a(n10264) );
no02f01  g4779 ( .o(n10267), .a(n10266), .b(n7340) );
oa12f01  g4780 ( .o(n10268), .a(n6148), .b(n10267), .c(n10265) );
ao12f01  g4781 ( .o(n10269), .a(n6131_1), .b(n6147), .c(_net_9377) );
na02f01  g4782 ( .o(n2965), .a(n10269), .b(n10268) );
in01f01  g4783 ( .o(n10271), .a(net_9508) );
ao22f01  g4784 ( .o(n10272), .a(n5743), .b(x1547), .c(n5742), .d(_net_9417) );
oa12f01  g4785 ( .o(n2970), .a(n10272), .b(n5741), .c(n10271) );
oa22f01  g4786 ( .o(n2975), .a(n7367), .b(n6720), .c(n7365_1), .d(n5537_1) );
ao12f01  g4787 ( .o(n10275), .a(n5658), .b(n5774), .c(x3949) );
oa12f01  g4788 ( .o(n2980), .a(n10275), .b(n5770), .c(n8931) );
oa22f01  g4789 ( .o(n2985), .a(n7756), .b(n6362), .c(n7755), .d(n9237) );
in01f01  g4790 ( .o(n10278), .a(_net_10206) );
ao12f01  g4791 ( .o(n10279), .a(n5658), .b(n6887), .c(x5722) );
oa12f01  g4792 ( .o(n2990), .a(n10279), .b(n6885_1), .c(n10278) );
in01f01  g4793 ( .o(n10281), .a(net_9952) );
in01f01  g4794 ( .o(n10282), .a(_net_234) );
oa22f01  g4795 ( .o(n2995), .a(n8831), .b(n10282), .c(n8829_1), .d(n10281) );
na02f01  g4796 ( .o(n10284), .a(n6056), .b(net_256) );
na02f01  g4797 ( .o(n10285), .a(n6055), .b(net_9984) );
ao22f01  g4798 ( .o(n10286), .a(n6062_1), .b(x4359), .c(n6060), .d(_net_10435) );
na04f01  g4799 ( .o(n3000), .a(n10286), .b(n10285), .c(n10284), .d(n6058) );
ao22f01  g4800 ( .o(n10288), .a(n5842), .b(net_9686), .c(n5841), .d(_net_124) );
na02f01  g4801 ( .o(n10289), .a(n5847), .b(net_9983) );
ao22f01  g4802 ( .o(n10290), .a(n5850), .b(net_9785), .c(n5849_1), .d(net_9884) );
na03f01  g4803 ( .o(n3005), .a(n10290), .b(n10289), .c(n10288) );
in01f01  g4804 ( .o(n10292), .a(net_10024) );
na03f01  g4805 ( .o(n10293), .a(n10292), .b(n7412), .c(n7396) );
in01f01  g4806 ( .o(n10294), .a(net_10023) );
na04f01  g4807 ( .o(n10295), .a(n10294), .b(n7399), .c(n7372), .d(n5897) );
na04f01  g4808 ( .o(n10296), .a(n7871_1), .b(n7389_1), .c(n7382), .d(n7379_1) );
no03f01  g4809 ( .o(n10297), .a(n10296), .b(n10295), .c(n10293) );
in01f01  g4810 ( .o(n10298), .a(_net_10463) );
no02f01  g4811 ( .o(n10299), .a(n10298), .b(_net_10033) );
no02f01  g4812 ( .o(n10300), .a(_net_10463), .b(n7372) );
in01f01  g4813 ( .o(n10301), .a(n10300) );
no02f01  g4814 ( .o(n10302), .a(n7382), .b(_net_10462) );
no02f01  g4815 ( .o(n10303), .a(n9719), .b(n9718) );
no02f01  g4816 ( .o(n10304), .a(n9719), .b(n9702) );
no02f01  g4817 ( .o(n10305), .a(_net_10032), .b(n9037) );
no02f01  g4818 ( .o(n10306), .a(n10305), .b(n9720) );
ao12f01  g4819 ( .o(n10307), .a(n10306), .b(n10302), .c(_net_10032) );
no02f01  g4820 ( .o(n10308), .a(n10307), .b(n10304) );
in01f01  g4821 ( .o(n10309), .a(n10308) );
no02f01  g4822 ( .o(n10310), .a(n10309), .b(n10303) );
na02f01  g4823 ( .o(n10311), .a(n10307), .b(_net_10462) );
oa12f01  g4824 ( .o(n10312), .a(n10311), .b(n10310), .c(n10302) );
ao12f01  g4825 ( .o(n10313), .a(n10299), .b(n10312), .c(n10301) );
na02f01  g4826 ( .o(n10314), .a(n10313), .b(n9048) );
no02f01  g4827 ( .o(n10315), .a(n10314), .b(_net_10465) );
ao12f01  g4828 ( .o(n3010), .a(n10297), .b(n10315), .c(n9054) );
na02f01  g4829 ( .o(n10317), .a(n6056), .b(net_242) );
na02f01  g4830 ( .o(n10318), .a(n6055), .b(net_9970) );
ao22f01  g4831 ( .o(n10319), .a(n6062_1), .b(x5427), .c(n6060), .d(_net_10421) );
na04f01  g4832 ( .o(n3015), .a(n10319), .b(n10318), .c(n10317), .d(n6058) );
in01f01  g4833 ( .o(n10321), .a(net_9251) );
na02f01  g4834 ( .o(n10322), .a(n6349), .b(x6599) );
na02f01  g4835 ( .o(n10323), .a(n6351_1), .b(x6599) );
oa22f01  g4836 ( .o(n3020), .a(n10323), .b(n10321), .c(n10322), .d(n6075) );
no02f01  g4837 ( .o(n10325), .a(n7240_1), .b(_net_9362) );
in01f01  g4838 ( .o(n10326), .a(_net_9362) );
no02f01  g4839 ( .o(n10327), .a(n7173_1), .b(n10326) );
no02f01  g4840 ( .o(n10328), .a(n10327), .b(n10325) );
no02f01  g4841 ( .o(n10329), .a(n10328), .b(n10257) );
na02f01  g4842 ( .o(n10330), .a(n10328), .b(n10257) );
na02f01  g4843 ( .o(n10331), .a(n10330), .b(n6148) );
ao12f01  g4844 ( .o(n10332), .a(n6131_1), .b(n6147), .c(_net_9370) );
oa12f01  g4845 ( .o(n3025), .a(n10332), .b(n10331), .c(n10329) );
ao12f01  g4846 ( .o(n10334), .a(n5658), .b(n5774), .c(x4117) );
oa12f01  g4847 ( .o(n3030), .a(n10334), .b(n5770), .c(n6994) );
na02f01  g4848 ( .o(n10336), .a(n7678), .b(_net_10439) );
na02f01  g4849 ( .o(n3043), .a(n10336), .b(n9318) );
no02f01  g4850 ( .o(n10338), .a(_net_9321), .b(_net_9320) );
no02f01  g4851 ( .o(n10339), .a(n8763), .b(n8332) );
no02f01  g4852 ( .o(n10340), .a(n10339), .b(n10338) );
no02f01  g4853 ( .o(n10341), .a(net_9157), .b(net_9158) );
in01f01  g4854 ( .o(n10342), .a(net_9157) );
no02f01  g4855 ( .o(n10343), .a(n10342), .b(n8643) );
no02f01  g4856 ( .o(n10344), .a(n10343), .b(n10341) );
na02f01  g4857 ( .o(n10345), .a(n10344), .b(n10340) );
in01f01  g4858 ( .o(n10346), .a(n10340) );
in01f01  g4859 ( .o(n10347), .a(n10344) );
na02f01  g4860 ( .o(n10348), .a(n10347), .b(n10346) );
na03f01  g4861 ( .o(n10349), .a(n10348), .b(n10345), .c(n8638) );
ao12f01  g4862 ( .o(n10350), .a(n7883), .b(n8637), .c(_net_9314) );
na02f01  g4863 ( .o(n3048), .a(n10350), .b(n10349) );
in01f01  g4864 ( .o(n10352), .a(_net_10414) );
ao12f01  g4865 ( .o(n10353), .a(n5658), .b(n6052_1), .c(x5850) );
oa12f01  g4866 ( .o(n3053), .a(n10353), .b(n6048), .c(n10352) );
na03f01  g4867 ( .o(n10355), .a(n5880), .b(n5879), .c(net_9533) );
in01f01  g4868 ( .o(n10356), .a(n5859) );
no02f01  g4869 ( .o(n10357), .a(n10356), .b(n5889) );
ao12f01  g4870 ( .o(n10358), .a(_net_9250), .b(n5889), .c(n5489) );
ao22f01  g4871 ( .o(n10359), .a(n10358), .b(n5865), .c(n10357), .d(n5857) );
na03f01  g4872 ( .o(n10360), .a(n5892), .b(n8399_1), .c(net_9533) );
oa12f01  g4873 ( .o(n10361), .a(n5871), .b(n8411), .c(_net_9250) );
na03f01  g4874 ( .o(n10362), .a(n10361), .b(net_9533), .c(n5489) );
na04f01  g4875 ( .o(n3058), .a(n10362), .b(n10360), .c(n10359), .d(n10355) );
in01f01  g4876 ( .o(n10364), .a(net_221) );
in01f01  g4877 ( .o(n10365), .a(net_9271) );
na02f01  g4878 ( .o(n10366), .a(n10365), .b(_net_9272) );
na03f01  g4879 ( .o(n10367), .a(n10366), .b(net_9271), .c(x6599) );
in01f01  g4880 ( .o(n10368), .a(net_220) );
no02f01  g4881 ( .o(n10369), .a(n10368), .b(n10364) );
in01f01  g4882 ( .o(n10370), .a(n10369) );
na02f01  g4883 ( .o(n10371), .a(n10368), .b(n10364) );
na02f01  g4884 ( .o(n10372), .a(n10371), .b(n10370) );
na03f01  g4885 ( .o(n10373), .a(n10365), .b(n7754), .c(x6599) );
oa22f01  g4886 ( .o(n3063), .a(n10373), .b(n10364), .c(n10372), .d(n10367) );
no02f01  g4887 ( .o(n10375), .a(n7763_1), .b(n8661) );
no02f01  g4888 ( .o(n10376), .a(_net_10160), .b(_net_9736) );
in01f01  g4889 ( .o(n10377), .a(n10376) );
no02f01  g4890 ( .o(n10378), .a(_net_9735), .b(_net_10159) );
in01f01  g4891 ( .o(n10379), .a(_net_9735) );
no02f01  g4892 ( .o(n10380), .a(n10379), .b(n7765) );
na02f01  g4893 ( .o(n10381), .a(n10379), .b(n7765) );
oa12f01  g4894 ( .o(n10382), .a(n10381), .b(n10380), .c(n8533) );
no04f01  g4895 ( .o(n10383), .a(n8534_1), .b(n8523), .c(n8135_1), .d(n8133) );
in01f01  g4896 ( .o(n10384), .a(n8534_1) );
na02f01  g4897 ( .o(n10385), .a(n10384), .b(n8528) );
na02f01  g4898 ( .o(n10386), .a(n10382), .b(n10385) );
no02f01  g4899 ( .o(n10387), .a(n10386), .b(n10383) );
oa22f01  g4900 ( .o(n10388), .a(n10387), .b(n10378), .c(n10382), .d(n7765) );
ao12f01  g4901 ( .o(n10389), .a(n10375), .b(n10388), .c(n10377) );
no02f01  g4902 ( .o(n10390), .a(n10389), .b(n7820) );
na02f01  g4903 ( .o(n10391), .a(n10390), .b(_net_10162) );
ao12f01  g4904 ( .o(n10392), .a(n6746), .b(n10391), .c(n9658) );
oa12f01  g4905 ( .o(n10393), .a(n10392), .b(n10391), .c(n9658) );
no02f01  g4906 ( .o(n10394), .a(n8541), .b(_net_10159) );
na02f01  g4907 ( .o(n10395), .a(n10394), .b(n7763_1) );
no02f01  g4908 ( .o(n10396), .a(n10395), .b(_net_10161) );
na03f01  g4909 ( .o(n10397), .a(n10396), .b(n9361), .c(_net_10163) );
in01f01  g4910 ( .o(n10398), .a(n6750) );
ao12f01  g4911 ( .o(n10399), .a(_net_10163), .b(n10396), .c(n9361) );
no02f01  g4912 ( .o(n10400), .a(n10399), .b(n10398) );
ao22f01  g4913 ( .o(n10401), .a(n10400), .b(n10397), .c(n6760), .d(_net_10163) );
na02f01  g4914 ( .o(n3068), .a(n10401), .b(n10393) );
na02f01  g4915 ( .o(n10403), .a(n8200_1), .b(n7029) );
na02f01  g4916 ( .o(n10404), .a(n5707), .b(n7029) );
na03f01  g4917 ( .o(n10405), .a(n10404), .b(n8183), .c(n9931) );
na02f01  g4918 ( .o(n10406), .a(n8202), .b(_net_10362) );
na03f01  g4919 ( .o(n3077), .a(n10406), .b(n10405), .c(n10403) );
ao12f01  g4920 ( .o(n10408), .a(n5658), .b(n7844), .c(_net_254) );
ao22f01  g4921 ( .o(n10409), .a(n7847), .b(x4520), .c(n7846), .d(net_9816) );
na02f01  g4922 ( .o(n3082), .a(n10409), .b(n10408) );
in01f01  g4923 ( .o(n10411), .a(_net_10309) );
ao12f01  g4924 ( .o(n10412), .a(n5658), .b(n5774), .c(x5850) );
oa12f01  g4925 ( .o(n3087), .a(n10412), .b(n5770), .c(n10411) );
in01f01  g4926 ( .o(n10414), .a(_net_10107) );
ao12f01  g4927 ( .o(n10415), .a(n5658), .b(n6160_1), .c(x5364) );
oa12f01  g4928 ( .o(n3092), .a(n10415), .b(n6159), .c(n10414) );
na02f01  g4929 ( .o(n10417), .a(n7353), .b(x5427) );
na02f01  g4930 ( .o(n10418), .a(n7352), .b(net_9673) );
ao22f01  g4931 ( .o(n10419), .a(n7358), .b(net_242), .c(n7357), .d(_net_10106) );
na04f01  g4932 ( .o(n3101), .a(n10419), .b(n10418), .c(n10417), .d(n7355_1) );
no03f01  g4933 ( .o(n10421), .a(_net_9248), .b(_net_9247), .c(_net_9249) );
in01f01  g4934 ( .o(n10422), .a(n10421) );
no02f01  g4935 ( .o(n10423), .a(n10422), .b(n10128) );
in01f01  g4936 ( .o(n10424), .a(_net_9235) );
no04f01  g4937 ( .o(n10425), .a(n10131), .b(n8451), .c(n10424), .d(_net_9236) );
no02f01  g4938 ( .o(n10426), .a(n6495), .b(n6491) );
no04f01  g4939 ( .o(n10427), .a(n10426), .b(n8453), .c(n8450), .d(_net_9235) );
oa12f01  g4940 ( .o(n10428), .a(n10423), .b(n10427), .c(n10425) );
oa12f01  g4941 ( .o(n3106), .a(n6682), .b(n10428), .c(_net_9238) );
na04f01  g4942 ( .o(n10430), .a(n8021_1), .b(n8017), .c(n8028), .d(n1521) );
no02f01  g4943 ( .o(n10431), .a(net_9184), .b(net_9182) );
in01f01  g4944 ( .o(n10432), .a(n10431) );
no02f01  g4945 ( .o(n10433), .a(net_9184), .b(_net_9183) );
ao12f01  g4946 ( .o(n10434), .a(n10433), .b(n10431), .c(n8025) );
oa12f01  g4947 ( .o(n10435), .a(n10434), .b(n10432), .c(n10430) );
no02f01  g4948 ( .o(n3111), .a(n10435), .b(n7701) );
no02f01  g4949 ( .o(n10437), .a(n9810), .b(_net_9294) );
na02f01  g4950 ( .o(n10438), .a(n9813), .b(n8809_1) );
oa22f01  g4951 ( .o(n3116), .a(n10438), .b(n10437), .c(n8817), .d(n7605_1) );
no02f01  g4952 ( .o(n3121), .a(net_9650), .b(net_9151) );
ao12f01  g4953 ( .o(n10441), .a(n7883), .b(n7923), .c(_net_9315) );
oa12f01  g4954 ( .o(n3126), .a(n10441), .b(n7925_1), .c(n8759) );
na03f01  g4955 ( .o(n10443), .a(net_9277), .b(net_9276), .c(net_9278) );
no03f01  g4956 ( .o(n3131), .a(n10443), .b(net_9275), .c(net_9274) );
oa22f01  g4957 ( .o(n3136), .a(n5907), .b(n7399), .c(n5905), .d(n5621) );
no02f01  g4958 ( .o(n10446), .a(n9820), .b(n8810) );
oa12f01  g4959 ( .o(n10447), .a(n10446), .b(n9818), .c(_net_9298) );
oa12f01  g4960 ( .o(n3151), .a(n10447), .b(n8817), .c(n7536) );
ao12f01  g4961 ( .o(n10449), .a(n5658), .b(n5678), .c(net_260) );
ao22f01  g4962 ( .o(n10450), .a(n5681_1), .b(x4041), .c(n5680), .d(net_9723) );
na02f01  g4963 ( .o(n3156), .a(n10450), .b(n10449) );
na02f01  g4964 ( .o(n10452), .a(n6056), .b(net_235) );
na02f01  g4965 ( .o(n10453), .a(n6055), .b(net_9963) );
ao22f01  g4966 ( .o(n10454), .a(n6062_1), .b(x5850), .c(n6060), .d(_net_10414) );
na04f01  g4967 ( .o(n3166), .a(n10454), .b(n10453), .c(n10452), .d(n6058) );
na02f01  g4968 ( .o(n10456), .a(n5749), .b(_net_10117) );
na02f01  g4969 ( .o(n3171), .a(n10456), .b(n5751) );
ao22f01  g4970 ( .o(n10458), .a(n5842), .b(net_9712), .c(n5841), .d(_net_152) );
na02f01  g4971 ( .o(n10459), .a(n5847), .b(net_10009) );
ao22f01  g4972 ( .o(n10460), .a(n5850), .b(net_9811), .c(n5849_1), .d(net_9910) );
na03f01  g4973 ( .o(n3176), .a(n10460), .b(n10459), .c(n10458) );
in01f01  g4974 ( .o(n10462), .a(net_10068) );
in01f01  g4975 ( .o(n10463), .a(_net_9660) );
na02f01  g4976 ( .o(n10464), .a(net_9659), .b(n10463) );
ao12f01  g4977 ( .o(n3181), .a(n6155_1), .b(n10464), .c(n10462) );
no02f01  g4978 ( .o(n10466), .a(n8334), .b(n7882) );
no02f01  g4979 ( .o(n10467), .a(_net_9326), .b(_net_9325) );
no02f01  g4980 ( .o(n10468), .a(n10467), .b(n10466) );
no02f01  g4981 ( .o(n10469), .a(net_9152), .b(n9375) );
no02f01  g4982 ( .o(n10470), .a(n8339_1), .b(net_9153) );
no02f01  g4983 ( .o(n10471), .a(n10470), .b(n10469) );
in01f01  g4984 ( .o(n10472), .a(n10471) );
no02f01  g4985 ( .o(n10473), .a(n10472), .b(_net_9311) );
in01f01  g4986 ( .o(n10474), .a(n10473) );
na02f01  g4987 ( .o(n10475), .a(n10472), .b(_net_9311) );
na03f01  g4988 ( .o(n10476), .a(n10475), .b(n10474), .c(n10468) );
in01f01  g4989 ( .o(n10477), .a(n10468) );
in01f01  g4990 ( .o(n10478), .a(n10475) );
oa12f01  g4991 ( .o(n10479), .a(n10477), .b(n10478), .c(n10473) );
na03f01  g4992 ( .o(n10480), .a(n10479), .b(n10476), .c(n8638) );
ao12f01  g4993 ( .o(n10481), .a(n7883), .b(n8637), .c(_net_9319) );
na02f01  g4994 ( .o(n3186), .a(n10481), .b(n10480) );
no02f01  g4995 ( .o(n10483), .a(n6655), .b(n6611) );
in01f01  g4996 ( .o(n10484), .a(n10483) );
na02f01  g4997 ( .o(n10485), .a(n10484), .b(n6663) );
na02f01  g4998 ( .o(n10486), .a(n10483), .b(n6653) );
na02f01  g4999 ( .o(n3191), .a(n10486), .b(n10485) );
na02f01  g5000 ( .o(n10488), .a(n7937), .b(net_243) );
na02f01  g5001 ( .o(n10489), .a(n7936), .b(net_9773) );
ao22f01  g5002 ( .o(n10490), .a(n7943), .b(_net_10212), .c(n7942), .d(x5364) );
na04f01  g5003 ( .o(n3195), .a(n10490), .b(n10489), .c(n10488), .d(n7939) );
in01f01  g5004 ( .o(n10492), .a(net_10189) );
no04f01  g5005 ( .o(n10493), .a(_net_9644), .b(_net_9646), .c(_net_9645), .d(_net_9643) );
in01f01  g5006 ( .o(n10494), .a(n10493) );
no03f01  g5007 ( .o(n10495), .a(n8753), .b(_net_9642), .c(_net_9640) );
no02f01  g5008 ( .o(n10496), .a(_net_9638), .b(_net_9639) );
na04f01  g5009 ( .o(n10497), .a(n10496), .b(n10495), .c(n8744), .d(_net_9649) );
no03f01  g5010 ( .o(n10498), .a(n9492), .b(n8772_1), .c(_net_9637) );
na04f01  g5011 ( .o(n10499), .a(n10498), .b(n10496), .c(n8753), .d(n9786) );
ao12f01  g5012 ( .o(n10500), .a(n10494), .b(n10499), .c(n10497) );
na02f01  g5013 ( .o(n10501), .a(n10500), .b(net_10175) );
ao12f01  g5014 ( .o(n3200), .a(n8577_1), .b(n10501), .c(n10492) );
ao12f01  g5015 ( .o(n10503), .a(n5658), .b(n7844), .c(net_242) );
ao22f01  g5016 ( .o(n10504), .a(n7847), .b(x5427), .c(n7846), .d(net_9804) );
na02f01  g5017 ( .o(n3205), .a(n10504), .b(n10503) );
ao12f01  g5018 ( .o(n10506), .a(n5658), .b(n7844), .c(net_257) );
ao22f01  g5019 ( .o(n10507), .a(n7847), .b(x4285), .c(n7846), .d(net_9819) );
na02f01  g5020 ( .o(n3215), .a(n10507), .b(n10506) );
in01f01  g5021 ( .o(n10509), .a(net_9225) );
no03f01  g5022 ( .o(n10510), .a(n9919), .b(n10509), .c(n9918) );
oa12f01  g5023 ( .o(n10511), .a(n9903), .b(n10510), .c(net_9226) );
ao12f01  g5024 ( .o(n3225), .a(n10511), .b(n10510), .c(net_9226) );
ao12f01  g5025 ( .o(n10513), .a(n5658), .b(n6875_1), .c(_net_254) );
ao22f01  g5026 ( .o(n10514), .a(n6878), .b(x4520), .c(n6877), .d(net_9915) );
na02f01  g5027 ( .o(n3230), .a(n10514), .b(n10513) );
na02f01  g5028 ( .o(n10516), .a(n6038), .b(net_257) );
na02f01  g5029 ( .o(n10517), .a(n6037_1), .b(net_9886) );
ao22f01  g5030 ( .o(n10518), .a(n6044), .b(x4285), .c(n6042_1), .d(_net_10331) );
na04f01  g5031 ( .o(n3238), .a(n10518), .b(n10517), .c(n10516), .d(n6040) );
in01f01  g5032 ( .o(n10520), .a(net_10073) );
oa22f01  g5033 ( .o(n3243), .a(n6989_1), .b(n5513_1), .c(n6988), .d(n10520) );
in01f01  g5034 ( .o(n10522), .a(net_9656) );
na02f01  g5035 ( .o(n10523), .a(n8705), .b(net_9655) );
no02f01  g5036 ( .o(n10524), .a(n10523), .b(n10522) );
in01f01  g5037 ( .o(n10525), .a(n10523) );
no02f01  g5038 ( .o(n10526), .a(n10525), .b(net_9656) );
no03f01  g5039 ( .o(n3252), .a(n10526), .b(n10524), .c(net_9151) );
na02f01  g5040 ( .o(n10528), .a(_net_9299), .b(_net_176) );
na02f01  g5041 ( .o(n10529), .a(n7529_1), .b(n5990) );
no02f01  g5042 ( .o(n10530), .a(n7573), .b(n7571_1) );
no02f01  g5043 ( .o(n10531), .a(_net_169), .b(_net_9292) );
no02f01  g5044 ( .o(n10532), .a(n5983_1), .b(n7516) );
no02f01  g5045 ( .o(n10533), .a(_net_177), .b(_net_9300) );
oa22f01  g5046 ( .o(n10534), .a(n10533), .b(n10532), .c(n10531), .d(n10530) );
ao12f01  g5047 ( .o(n10535), .a(n10534), .b(n10529), .c(n10528) );
na02f01  g5048 ( .o(n10536), .a(n8473), .b(n8467_1) );
no02f01  g5049 ( .o(n10537), .a(n5916), .b(n6025) );
no02f01  g5050 ( .o(n10538), .a(_net_168), .b(_net_9291) );
no02f01  g5051 ( .o(n10539), .a(n7593), .b(n7592) );
no02f01  g5052 ( .o(n10540), .a(_net_9290), .b(_net_167) );
oa22f01  g5053 ( .o(n10541), .a(n10540), .b(n10539), .c(n10538), .d(n10537) );
in01f01  g5054 ( .o(n10542), .a(n8463) );
na02f01  g5055 ( .o(n10543), .a(n8477_1), .b(n8476) );
no03f01  g5056 ( .o(n10544), .a(n10543), .b(n8487), .c(n8481) );
na04f01  g5057 ( .o(n10545), .a(n10544), .b(n8471), .c(n10542), .d(n8457_1) );
no03f01  g5058 ( .o(n10546), .a(n10545), .b(n10541), .c(n10536) );
na02f01  g5059 ( .o(n10547), .a(n5924), .b(_net_9646) );
ao12f01  g5060 ( .o(n3257), .a(n10547), .b(n10546), .c(n10535) );
in01f01  g5061 ( .o(n10549), .a(_net_9192) );
oa22f01  g5062 ( .o(n3262), .a(n8349_1), .b(n8034), .c(n8347), .d(n10549) );
ao12f01  g5063 ( .o(n10551), .a(n5658), .b(n6875_1), .c(_net_261) );
ao22f01  g5064 ( .o(n10552), .a(n6878), .b(x3949), .c(n6877), .d(net_9922) );
na02f01  g5065 ( .o(n3267), .a(n10552), .b(n10551) );
na02f01  g5066 ( .o(n10554), .a(n7489), .b(n6514) );
oa12f01  g5067 ( .o(n4966), .a(n10554), .b(n10062), .c(n6514) );
oa12f01  g5068 ( .o(n10556), .a(x6599), .b(n4966), .c(net_9197) );
na02f01  g5069 ( .o(n10557), .a(n4966), .b(net_9197) );
ao12f01  g5070 ( .o(n3272), .a(n10556), .b(n10557), .c(n6515) );
na02f01  g5071 ( .o(n10559), .a(net_113), .b(_net_9606) );
in01f01  g5072 ( .o(n10560), .a(n7511) );
oa12f01  g5073 ( .o(n10561), .a(n10560), .b(n7624), .c(n7541) );
no02f01  g5074 ( .o(n10562), .a(n7505), .b(n7503) );
ao12f01  g5075 ( .o(n10563), .a(n10562), .b(n10561), .c(n7509_1) );
in01f01  g5076 ( .o(n10564), .a(n7541) );
ao12f01  g5077 ( .o(n10565), .a(n7511), .b(n7636_1), .c(n10564) );
in01f01  g5078 ( .o(n10566), .a(n10562) );
no03f01  g5079 ( .o(n10567), .a(n10566), .b(n10565), .c(n7508) );
oa12f01  g5080 ( .o(n10568), .a(n7500), .b(n10567), .c(n10563) );
na02f01  g5081 ( .o(n3277), .a(n10568), .b(n10559) );
na02f01  g5082 ( .o(n10570), .a(n6168), .b(_net_10247) );
na02f01  g5083 ( .o(n10571), .a(n6831_1), .b(n6781) );
na03f01  g5084 ( .o(n10572), .a(n10571), .b(n6833), .c(n6175) );
no02f01  g5085 ( .o(n10573), .a(n6786_1), .b(n6782_1) );
in01f01  g5086 ( .o(n10574), .a(n10573) );
na02f01  g5087 ( .o(n10575), .a(n10574), .b(n6792) );
oa12f01  g5088 ( .o(n10576), .a(n10573), .b(n6791_1), .c(n6788) );
na03f01  g5089 ( .o(n10577), .a(n10576), .b(n10575), .c(n6177_1) );
na03f01  g5090 ( .o(n3282), .a(n10577), .b(n10572), .c(n10570) );
ao22f01  g5091 ( .o(n10579), .a(n5842), .b(net_9663), .c(n5841), .d(net_101) );
na02f01  g5092 ( .o(n10580), .a(n5847), .b(net_9960) );
ao22f01  g5093 ( .o(n10581), .a(n5850), .b(net_9762), .c(n5849_1), .d(net_9861) );
na03f01  g5094 ( .o(n3287), .a(n10581), .b(n10580), .c(n10579) );
in01f01  g5095 ( .o(n10583), .a(_net_9193) );
in01f01  g5096 ( .o(n10584), .a(net_9184) );
oa22f01  g5097 ( .o(n3296), .a(n8349_1), .b(n10584), .c(n8347), .d(n10583) );
ao12f01  g5098 ( .o(n10586), .a(n5658), .b(n6887), .c(x4041) );
oa12f01  g5099 ( .o(n3305), .a(n10586), .b(n6885_1), .c(n9180) );
in01f01  g5100 ( .o(n10588), .a(net_10296) );
na02f01  g5101 ( .o(n10589), .a(net_10280), .b(net_264) );
ao12f01  g5102 ( .o(n3315), .a(n5911), .b(n10589), .c(n10588) );
oa22f01  g5103 ( .o(n3320), .a(n7367), .b(n5782_1), .c(n7365_1), .d(n5612) );
ao12f01  g5104 ( .o(n10592), .a(n5658), .b(n6875_1), .c(net_250) );
ao22f01  g5105 ( .o(n10593), .a(n6878), .b(x4851), .c(n6877), .d(net_9911) );
na02f01  g5106 ( .o(n3325), .a(n10593), .b(n10592) );
in01f01  g5107 ( .o(n10595), .a(n9197) );
no03f01  g5108 ( .o(n10596), .a(n9206), .b(n9203), .c(n10595) );
no02f01  g5109 ( .o(n10597), .a(n9207), .b(n9187) );
na02f01  g5110 ( .o(n10598), .a(n10597), .b(n10596) );
in01f01  g5111 ( .o(n10599), .a(n10596) );
in01f01  g5112 ( .o(n10600), .a(n10597) );
na02f01  g5113 ( .o(n10601), .a(n10600), .b(n10599) );
na02f01  g5114 ( .o(n3330), .a(n10601), .b(n10598) );
no03f01  g5115 ( .o(n10603), .a(n6474_1), .b(n8446), .c(n6463) );
no02f01  g5116 ( .o(n10604), .a(n6502), .b(n8446) );
na02f01  g5117 ( .o(n10605), .a(n10604), .b(n6508) );
oa12f01  g5118 ( .o(n10606), .a(n10604), .b(n6506), .c(_net_9248) );
na02f01  g5119 ( .o(n10607), .a(n10606), .b(n10605) );
no03f01  g5120 ( .o(n10608), .a(n7482), .b(n6485), .c(n8446) );
na03f01  g5121 ( .o(n10609), .a(n6860), .b(_net_9242), .c(_net_9236) );
no03f01  g5122 ( .o(n10610), .a(_net_9209), .b(n6520), .c(n8446) );
no02f01  g5123 ( .o(n10611), .a(n6477), .b(n8446) );
no03f01  g5124 ( .o(n10612), .a(n10611), .b(n10610), .c(n6678) );
in01f01  g5125 ( .o(n10613), .a(n6498_1) );
na02f01  g5126 ( .o(n10614), .a(n10613), .b(n6495) );
oa12f01  g5127 ( .o(n10615), .a(_net_9242), .b(n10614), .c(n6494) );
na03f01  g5128 ( .o(n10616), .a(n10615), .b(n10612), .c(n10609) );
no04f01  g5129 ( .o(n10617), .a(n10616), .b(n10608), .c(n10607), .d(n10603) );
no02f01  g5130 ( .o(n3335), .a(n10617), .b(n6526_1) );
oa22f01  g5131 ( .o(n3340), .a(n9353), .b(n5640), .c(n9352), .d(n8301_1) );
na02f01  g5132 ( .o(n10620), .a(n7937), .b(net_262) );
na02f01  g5133 ( .o(n10621), .a(n7936), .b(net_9792) );
ao22f01  g5134 ( .o(n10622), .a(n7943), .b(_net_10231), .c(n7942), .d(x3889) );
na04f01  g5135 ( .o(n3345), .a(n10622), .b(n10621), .c(n10620), .d(n7939) );
na02f01  g5136 ( .o(n10624), .a(n7358), .b(net_249) );
na02f01  g5137 ( .o(n10625), .a(n7352), .b(net_9680) );
ao22f01  g5138 ( .o(n10626), .a(n7357), .b(_net_10113), .c(n7353), .d(x4937) );
na04f01  g5139 ( .o(n3350), .a(n10626), .b(n10625), .c(n10624), .d(n7355_1) );
in01f01  g5140 ( .o(n10628), .a(_net_10531) );
ao12f01  g5141 ( .o(n10629), .a(n8082), .b(n8074), .c(n5496) );
na04f01  g5142 ( .o(n10630), .a(n8076_1), .b(_net_10538), .c(n5500_1), .d(x6157) );
oa12f01  g5143 ( .o(n3355), .a(n10630), .b(n10629), .c(n10628) );
na03f01  g5144 ( .o(n10632), .a(n8079), .b(n6570), .c(_net_10529) );
no02f01  g5145 ( .o(n3369), .a(n10632), .b(n5901) );
ao22f01  g5146 ( .o(n10634), .a(n9018), .b(_net_10443), .c(_net_10444), .d(n9017) );
no02f01  g5147 ( .o(n10635), .a(_net_10442), .b(n9013) );
ao22f01  g5148 ( .o(n10636), .a(n9014), .b(_net_8839), .c(_net_10442), .d(n9013) );
oa12f01  g5149 ( .o(n10637), .a(n10634), .b(n10636), .c(n10635) );
in01f01  g5150 ( .o(n10638), .a(_net_10443) );
in01f01  g5151 ( .o(n10639), .a(_net_10444) );
ao12f01  g5152 ( .o(n10640), .a(n9018), .b(_net_10444), .c(n9017) );
ao22f01  g5153 ( .o(n10641), .a(n10640), .b(n10638), .c(n10639), .d(_net_10458) );
ao22f01  g5154 ( .o(n10642), .a(net_10447), .b(n9036), .c(n9037), .d(net_10448) );
ao22f01  g5155 ( .o(n10643), .a(n9025), .b(_net_10445), .c(n9024), .d(_net_10446) );
na02f01  g5156 ( .o(n10644), .a(n10643), .b(n10642) );
ao12f01  g5157 ( .o(n10645), .a(n10644), .b(n10641), .c(n10637) );
in01f01  g5158 ( .o(n10646), .a(net_10450) );
oa12f01  g5159 ( .o(n10647), .a(_net_10463), .b(_net_10464), .c(n10646) );
oa22f01  g5160 ( .o(n10648), .a(n10647), .b(net_10449), .c(n9048), .d(net_10450) );
in01f01  g5161 ( .o(n10649), .a(_net_10465) );
ao22f01  g5162 ( .o(n10650), .a(n9054), .b(_net_10452), .c(n10649), .d(_net_10451) );
in01f01  g5163 ( .o(n10651), .a(_net_10452) );
oa12f01  g5164 ( .o(n10652), .a(_net_10465), .b(_net_10466), .c(n10651) );
oa22f01  g5165 ( .o(n10653), .a(n10652), .b(_net_10451), .c(n9054), .d(_net_10452) );
ao12f01  g5166 ( .o(n10654), .a(n10653), .b(n10650), .c(n10648) );
in01f01  g5167 ( .o(n10655), .a(_net_10446) );
oa12f01  g5168 ( .o(n10656), .a(_net_10459), .b(_net_10460), .c(n10655) );
oa22f01  g5169 ( .o(n10657), .a(n10656), .b(_net_10445), .c(n9024), .d(_net_10446) );
in01f01  g5170 ( .o(n10658), .a(net_10448) );
oa12f01  g5171 ( .o(n10659), .a(_net_10461), .b(_net_10462), .c(n10658) );
oa22f01  g5172 ( .o(n10660), .a(n10659), .b(net_10447), .c(n9037), .d(net_10448) );
ao12f01  g5173 ( .o(n10661), .a(n10660), .b(n10657), .c(n10642) );
na02f01  g5174 ( .o(n10662), .a(n10661), .b(n10654) );
in01f01  g5175 ( .o(n10663), .a(n10650) );
in01f01  g5176 ( .o(n10664), .a(net_10449) );
oa22f01  g5177 ( .o(n10665), .a(n10664), .b(_net_10463), .c(_net_10464), .d(n10646) );
oa12f01  g5178 ( .o(n10666), .a(n10654), .b(n10665), .c(n10663) );
oa12f01  g5179 ( .o(n3374), .a(n10666), .b(n10662), .c(n10645) );
no02f01  g5180 ( .o(n10668), .a(n7215), .b(n7140) );
no02f01  g5181 ( .o(n10669), .a(n7192_1), .b(n7139) );
no02f01  g5182 ( .o(n10670), .a(n10669), .b(n10668) );
no02f01  g5183 ( .o(n10671), .a(n10670), .b(n10239) );
na02f01  g5184 ( .o(n10672), .a(n10670), .b(n10239) );
na02f01  g5185 ( .o(n10673), .a(n10672), .b(n6148) );
ao12f01  g5186 ( .o(n10674), .a(n6131_1), .b(n6147), .c(net_9364) );
oa12f01  g5187 ( .o(n3379), .a(n10674), .b(n10673), .c(n10671) );
na02f01  g5188 ( .o(n10676), .a(n8881), .b(n8856) );
na02f01  g5189 ( .o(n10677), .a(n8891), .b(n10676) );
na02f01  g5190 ( .o(n10678), .a(n10677), .b(n8908) );
no02f01  g5191 ( .o(n10679), .a(n8913), .b(n8882) );
in01f01  g5192 ( .o(n10680), .a(n10679) );
na02f01  g5193 ( .o(n10681), .a(n10680), .b(n10678) );
na03f01  g5194 ( .o(n10682), .a(n10679), .b(n10677), .c(n8908) );
na02f01  g5195 ( .o(n3384), .a(n10682), .b(n10681) );
oa12f01  g5196 ( .o(n10684), .a(n8074), .b(n5497), .c(net_10533) );
in01f01  g5197 ( .o(n10685), .a(net_10533) );
no03f01  g5198 ( .o(n10686), .a(n8081_1), .b(n8077), .c(n10685) );
ao12f01  g5199 ( .o(n10687), .a(n10686), .b(net_10532), .c(x6599) );
na02f01  g5200 ( .o(n3389), .a(n10687), .b(n10684) );
oa22f01  g5201 ( .o(n3394), .a(n5694), .b(n5815_1), .c(n5692), .d(n5640) );
oa22f01  g5202 ( .o(n3399), .a(n5907), .b(n6588), .c(n5905), .d(n5576) );
ao12f01  g5203 ( .o(n10691), .a(n5658), .b(n6052_1), .c(x4449) );
oa12f01  g5204 ( .o(n3404), .a(n10691), .b(n6048), .c(n8209) );
in01f01  g5205 ( .o(n10693), .a(net_10066) );
in01f01  g5206 ( .o(n10694), .a(net_10070) );
oa22f01  g5207 ( .o(n10695), .a(n10694), .b(n6985_1), .c(n10693), .d(n8282) );
ao12f01  g5208 ( .o(n10696), .a(n10695), .b(net_10087), .c(net_10069) );
in01f01  g5209 ( .o(n10697), .a(net_10086) );
in01f01  g5210 ( .o(n10698), .a(net_10082) );
in01f01  g5211 ( .o(n10699), .a(net_10064) );
oa22f01  g5212 ( .o(n10700), .a(n10699), .b(n10698), .c(n10697), .d(n10462) );
in01f01  g5213 ( .o(n10701), .a(net_10067) );
in01f01  g5214 ( .o(n10702), .a(net_10085) );
oa22f01  g5215 ( .o(n10703), .a(n10702), .b(n10701), .c(n9238), .d(n6152) );
no02f01  g5216 ( .o(n10704), .a(n10703), .b(n10700) );
no04f01  g5217 ( .o(n10705), .a(_net_9958), .b(_net_10057), .c(net_9760), .d(net_9859) );
ao22f01  g5218 ( .o(n10706), .a(net_10071), .b(net_10089), .c(net_10063), .d(net_10081) );
na04f01  g5219 ( .o(n3409), .a(n10706), .b(n10705), .c(n10704), .d(n10696) );
in01f01  g5220 ( .o(n10708), .a(_net_10100) );
ao12f01  g5221 ( .o(n10709), .a(n5658), .b(n6160_1), .c(x5790) );
oa12f01  g5222 ( .o(n3421), .a(n10709), .b(n6159), .c(n10708) );
in01f01  g5223 ( .o(n10711), .a(net_10392) );
oa22f01  g5224 ( .o(n3430), .a(n10211), .b(n5576), .c(n10210), .d(n10711) );
in01f01  g5225 ( .o(n10713), .a(net_210) );
oa22f01  g5226 ( .o(n3435), .a(n7756), .b(n6355), .c(n7755), .d(n10713) );
na02f01  g5227 ( .o(n10715), .a(n6020), .b(n5998_1) );
oa12f01  g5228 ( .o(n4293), .a(n10715), .b(n6020), .c(n5989) );
na02f01  g5229 ( .o(n10717), .a(n4293), .b(n7991) );
no02f01  g5230 ( .o(n10718), .a(n9464), .b(net_9524) );
no02f01  g5231 ( .o(n10719), .a(n9620), .b(n9457) );
no03f01  g5232 ( .o(n10720), .a(n10719), .b(n10718), .c(n7999) );
oa12f01  g5233 ( .o(n10721), .a(x6599), .b(n8002), .c(n9457) );
no02f01  g5234 ( .o(n10722), .a(n10721), .b(n10720) );
na02f01  g5235 ( .o(n3445), .a(n10722), .b(n10717) );
ao12f01  g5236 ( .o(n10724), .a(n5658), .b(n6875_1), .c(_net_255) );
ao22f01  g5237 ( .o(n10725), .a(n6878), .b(x4449), .c(n6877), .d(net_9916) );
na02f01  g5238 ( .o(n3450), .a(n10725), .b(n10724) );
in01f01  g5239 ( .o(n10727), .a(n7045) );
na02f01  g5240 ( .o(n10728), .a(n10727), .b(n7038) );
no02f01  g5241 ( .o(n10729), .a(n7043), .b(n7011) );
in01f01  g5242 ( .o(n10730), .a(n10729) );
na02f01  g5243 ( .o(n10731), .a(n10730), .b(n10728) );
na03f01  g5244 ( .o(n10732), .a(n10729), .b(n10727), .c(n7038) );
na02f01  g5245 ( .o(n3460), .a(n10732), .b(n10731) );
na02f01  g5246 ( .o(n10734), .a(n7937), .b(net_256) );
na02f01  g5247 ( .o(n10735), .a(n7936), .b(net_9786) );
ao22f01  g5248 ( .o(n10736), .a(n7943), .b(_net_10225), .c(n7942), .d(x4359) );
na04f01  g5249 ( .o(n3470), .a(n10736), .b(n10735), .c(n10734), .d(n7939) );
in01f01  g5250 ( .o(n10738), .a(net_10387) );
oa22f01  g5251 ( .o(n3475), .a(n10211), .b(n5567_1), .c(n10210), .d(n10738) );
in01f01  g5252 ( .o(n3480), .a(_net_10324) );
in01f01  g5253 ( .o(n10741), .a(net_10499) );
oa22f01  g5254 ( .o(n3485), .a(n7467), .b(n5612), .c(n7465_1), .d(n10741) );
no02f01  g5255 ( .o(n7365), .a(n6021), .b(n8918) );
in01f01  g5256 ( .o(n10744), .a(n7365) );
no02f01  g5257 ( .o(n3490), .a(n10744), .b(n5927) );
no02f01  g5258 ( .o(n3499), .a(n8578), .b(_net_9606) );
oa22f01  g5259 ( .o(n3504), .a(n7480_1), .b(n5799), .c(n7478), .d(n5640) );
ao12f01  g5260 ( .o(n10748), .a(n5658), .b(n6532), .c(net_249) );
ao22f01  g5261 ( .o(n10749), .a(n6535), .b(x4937), .c(n6534), .d(net_10009) );
na02f01  g5262 ( .o(n3513), .a(n10749), .b(n10748) );
na02f01  g5263 ( .o(n10751), .a(n7937), .b(net_252) );
na02f01  g5264 ( .o(n10752), .a(n7936), .b(net_9782) );
ao22f01  g5265 ( .o(n10753), .a(n7943), .b(_net_10221), .c(n7942), .d(x4694) );
na04f01  g5266 ( .o(n3518), .a(n10753), .b(n10752), .c(n10751), .d(n7939) );
na02f01  g5267 ( .o(n10755), .a(n9399), .b(n8090) );
na02f01  g5268 ( .o(n10756), .a(n10755), .b(n9401) );
oa22f01  g5269 ( .o(n3523), .a(n10756), .b(n9397), .c(n9407), .d(n8090) );
in01f01  g5270 ( .o(n10758), .a(net_10496) );
oa22f01  g5271 ( .o(n3528), .a(n7467), .b(n5525), .c(n7465_1), .d(n10758) );
na02f01  g5272 ( .o(n10760), .a(n6020), .b(n6634_1) );
oa12f01  g5273 ( .o(n8621), .a(n10760), .b(n6020), .c(n8466) );
na02f01  g5274 ( .o(n10762), .a(n8621), .b(n7991) );
oa12f01  g5275 ( .o(n10763), .a(net_9522), .b(n9461), .c(_net_9521) );
ao12f01  g5276 ( .o(n10764), .a(n7999), .b(n10763), .c(n9463) );
oa12f01  g5277 ( .o(n10765), .a(x6599), .b(n8002), .c(n9458) );
no02f01  g5278 ( .o(n10766), .a(n10765), .b(n10764) );
na02f01  g5279 ( .o(n3533), .a(n10766), .b(n10762) );
na02f01  g5280 ( .o(n10768), .a(n7937), .b(_net_255) );
na02f01  g5281 ( .o(n10769), .a(n7936), .b(net_9785) );
ao22f01  g5282 ( .o(n10770), .a(n7943), .b(_net_10224), .c(n7942), .d(x4449) );
na04f01  g5283 ( .o(n3538), .a(n10770), .b(n10769), .c(n10768), .d(n7939) );
in01f01  g5284 ( .o(n10772), .a(_net_10218) );
ao12f01  g5285 ( .o(n10773), .a(n5658), .b(n6887), .c(x4937) );
oa12f01  g5286 ( .o(n3543), .a(n10773), .b(n6885_1), .c(n10772) );
na02f01  g5287 ( .o(n10775), .a(n6695), .b(n6691) );
na04f01  g5288 ( .o(n10776), .a(n7651), .b(n6689_1), .c(n7650_1), .d(n6671) );
ao12f01  g5289 ( .o(n10777), .a(n10776), .b(n10775), .c(_net_9204) );
no02f01  g5290 ( .o(n3548), .a(n10777), .b(n6686) );
in01f01  g5291 ( .o(n10779), .a(net_10195) );
na02f01  g5292 ( .o(n10780), .a(_net_9117), .b(net_10175) );
ao12f01  g5293 ( .o(n3553), .a(n8577_1), .b(n10780), .c(n10779) );
in01f01  g5294 ( .o(n10782), .a(net_10394) );
oa22f01  g5295 ( .o(n3558), .a(n10211), .b(n5612), .c(n10210), .d(n10782) );
oa12f01  g5296 ( .o(n10784), .a(_net_9641), .b(n9542), .c(n9495) );
no04f01  g5297 ( .o(n10785), .a(n8751), .b(n7975), .c(n7969), .d(n7964) );
oa12f01  g5298 ( .o(n10786), .a(n10785), .b(n8747_1), .c(_net_9641) );
no02f01  g5299 ( .o(n10787), .a(n9546), .b(n8753) );
ao22f01  g5300 ( .o(n10788), .a(n10787), .b(n8774), .c(n9496), .d(_net_9641) );
na03f01  g5301 ( .o(n10789), .a(n10788), .b(n10786), .c(n10784) );
na02f01  g5302 ( .o(n10790), .a(n10789), .b(x6599) );
no02f01  g5303 ( .o(n3563), .a(n10790), .b(n2827) );
ao12f01  g5304 ( .o(n10792), .a(n5658), .b(n6887), .c(x4359) );
oa12f01  g5305 ( .o(n3568), .a(n10792), .b(n6885_1), .c(n9205) );
in01f01  g5306 ( .o(n10794), .a(net_10284) );
oa22f01  g5307 ( .o(n3573), .a(n9353), .b(n5637), .c(n9352), .d(n10794) );
ao12f01  g5308 ( .o(n10796), .a(n5658), .b(n6160_1), .c(x3949) );
oa12f01  g5309 ( .o(n3578), .a(n10796), .b(n6159), .c(n6667) );
ao12f01  g5310 ( .o(n10798), .a(n5658), .b(n6887), .c(x4781) );
oa12f01  g5311 ( .o(n3583), .a(n10798), .b(n6885_1), .c(n8960) );
in01f01  g5312 ( .o(n10800), .a(net_10294) );
na02f01  g5313 ( .o(n10801), .a(n10500), .b(net_10280) );
ao12f01  g5314 ( .o(n3588), .a(n5911), .b(n10801), .c(n10800) );
ao22f01  g5315 ( .o(n10803), .a(n5842), .b(_net_9731), .c(n5841), .d(_net_172) );
na02f01  g5316 ( .o(n10804), .a(n5847), .b(_net_10028) );
ao22f01  g5317 ( .o(n10805), .a(n5850), .b(_net_9830), .c(n5849_1), .d(_net_9929) );
na03f01  g5318 ( .o(n3593), .a(n10805), .b(n10804), .c(n10803) );
in01f01  g5319 ( .o(n10807), .a(_net_10096) );
ao12f01  g5320 ( .o(n10808), .a(n5658), .b(n6160_1), .c(x6028) );
oa12f01  g5321 ( .o(n3598), .a(n10808), .b(n6159), .c(n10807) );
in01f01  g5322 ( .o(n10810), .a(net_9859) );
in01f01  g5323 ( .o(n10811), .a(net_9858) );
na02f01  g5324 ( .o(n3603), .a(n10811), .b(n10810) );
na02f01  g5325 ( .o(n10813), .a(n7358), .b(net_257) );
na02f01  g5326 ( .o(n10814), .a(n7352), .b(net_9688) );
ao22f01  g5327 ( .o(n10815), .a(n7357), .b(_net_10121), .c(n7353), .d(x4285) );
na04f01  g5328 ( .o(n3608), .a(n10815), .b(n10814), .c(n10813), .d(n7355_1) );
oa22f01  g5329 ( .o(n3613), .a(n7467), .b(n5640), .c(n7465_1), .d(n8298) );
in01f01  g5330 ( .o(n10818), .a(net_218) );
oa22f01  g5331 ( .o(n3618), .a(n7756), .b(n5787_1), .c(n7755), .d(n10818) );
ao12f01  g5332 ( .o(n10820), .a(n7606), .b(n6028_1), .c(n6617) );
oa12f01  g5333 ( .o(n3628), .a(n10820), .b(n6022), .c(n8468) );
in01f01  g5334 ( .o(n10822), .a(x715) );
na02f01  g5335 ( .o(n10823), .a(n10164), .b(n7097) );
oa12f01  g5336 ( .o(n10824), .a(n10823), .b(n10164), .c(net_9364) );
no02f01  g5337 ( .o(n10825), .a(n10173), .b(n10161) );
ao22f01  g5338 ( .o(n10826), .a(n10825), .b(n10824), .c(n10161), .d(n7234) );
na03f01  g5339 ( .o(n10827), .a(n10158), .b(n10155), .c(n10156) );
oa22f01  g5340 ( .o(n3638), .a(n10827), .b(n10826), .c(n10155), .d(n10822) );
oa22f01  g5341 ( .o(n3642), .a(n6989_1), .b(n5552_1), .c(n6988), .d(n10697) );
in01f01  g5342 ( .o(n10830), .a(_net_10313) );
ao12f01  g5343 ( .o(n10831), .a(n5658), .b(n5774), .c(x5601) );
oa12f01  g5344 ( .o(n3652), .a(n10831), .b(n5770), .c(n10830) );
in01f01  g5345 ( .o(n10833), .a(net_216) );
ao22f01  g5346 ( .o(n10834), .a(n8047), .b(net_10066), .c(n6564), .d(net_10088) );
oa12f01  g5347 ( .o(n10835), .a(n10834), .b(n6563), .c(n10833) );
na02f01  g5348 ( .o(n10836), .a(n6584_1), .b(net_9784) );
na02f01  g5349 ( .o(n10837), .a(n6602), .b(net_10014) );
ao22f01  g5350 ( .o(n10838), .a(n6606), .b(net_9946), .c(n6597), .d(net_9748) );
na03f01  g5351 ( .o(n10839), .a(n10838), .b(n10837), .c(n10836) );
no02f01  g5352 ( .o(n10840), .a(n10839), .b(n10835) );
ao22f01  g5353 ( .o(n10841), .a(n6585), .b(net_9717), .c(n6573), .d(net_9883) );
ao22f01  g5354 ( .o(n10842), .a(n6582), .b(net_9915), .c(n6555), .d(net_9982) );
in01f01  g5355 ( .o(n10843), .a(net_9816) );
oa22f01  g5356 ( .o(n10844), .a(n6591), .b(n8620), .c(n9978), .d(n10843) );
in01f01  g5357 ( .o(n10845), .a(net_9847) );
na02f01  g5358 ( .o(n10846), .a(n6577), .b(net_9685) );
oa12f01  g5359 ( .o(n10847), .a(n10846), .b(n6600), .c(n10845) );
no02f01  g5360 ( .o(n10848), .a(n10847), .b(n10844) );
na04f01  g5361 ( .o(n3657), .a(n10848), .b(n10842), .c(n10841), .d(n10840) );
na02f01  g5362 ( .o(n10850), .a(n8756), .b(_net_8824) );
ao12f01  g5363 ( .o(n3662), .a(n5658), .b(n10850), .c(n8637) );
ao12f01  g5364 ( .o(n10852), .a(n5658), .b(n6532), .c(net_256) );
ao22f01  g5365 ( .o(n10853), .a(n6535), .b(x4359), .c(n6534), .d(net_10016) );
na02f01  g5366 ( .o(n3667), .a(n10853), .b(n10852) );
na02f01  g5367 ( .o(n10855), .a(n7937), .b(net_245) );
na02f01  g5368 ( .o(n10856), .a(n7936), .b(net_9775) );
ao22f01  g5369 ( .o(n10857), .a(n7943), .b(_net_10214), .c(n7942), .d(x5225) );
na04f01  g5370 ( .o(n3672), .a(n10857), .b(n10856), .c(n10855), .d(n7939) );
na02f01  g5371 ( .o(n10859), .a(n7937), .b(net_239) );
na02f01  g5372 ( .o(n10860), .a(n7936), .b(net_9769) );
ao22f01  g5373 ( .o(n10861), .a(n7943), .b(_net_10208), .c(n7942), .d(x5601) );
na04f01  g5374 ( .o(n3677), .a(n10861), .b(n10860), .c(n10859), .d(n7939) );
no02f01  g5375 ( .o(n10863), .a(n9199), .b(n9195) );
in01f01  g5376 ( .o(n10864), .a(n10863) );
oa12f01  g5377 ( .o(n10865), .a(n10864), .b(n9201), .c(n9192) );
in01f01  g5378 ( .o(n10866), .a(n9192) );
in01f01  g5379 ( .o(n10867), .a(n9201) );
na03f01  g5380 ( .o(n10868), .a(n10863), .b(n10867), .c(n10866) );
na02f01  g5381 ( .o(n3682), .a(n10868), .b(n10865) );
no02f01  g5382 ( .o(n10870), .a(n7406), .b(n7405) );
ao12f01  g5383 ( .o(n10871), .a(n7418_1), .b(n10870), .c(n7411) );
in01f01  g5384 ( .o(n10872), .a(n10871) );
no02f01  g5385 ( .o(n10873), .a(n7381), .b(n7407) );
ao12f01  g5386 ( .o(n10874), .a(n7875), .b(n10873), .c(n10872) );
oa12f01  g5387 ( .o(n10875), .a(n10874), .b(n10873), .c(n10872) );
na02f01  g5388 ( .o(n10876), .a(n7441_1), .b(_net_10473) );
na02f01  g5389 ( .o(n10877), .a(n10876), .b(n7443) );
ao22f01  g5390 ( .o(n10878), .a(n10877), .b(n7450), .c(n7453), .d(_net_10473) );
na02f01  g5391 ( .o(n3687), .a(n10878), .b(n10875) );
no02f01  g5392 ( .o(n10880), .a(n8216), .b(n8214_1) );
in01f01  g5393 ( .o(n10881), .a(n10880) );
na02f01  g5394 ( .o(n10882), .a(n10881), .b(n8235_1) );
in01f01  g5395 ( .o(n10883), .a(n8235_1) );
na02f01  g5396 ( .o(n10884), .a(n10880), .b(n10883) );
na02f01  g5397 ( .o(n3692), .a(n10884), .b(n10882) );
oa22f01  g5398 ( .o(n3697), .a(n5694), .b(n9976), .c(n5692), .d(n5603) );
in01f01  g5399 ( .o(n10887), .a(_net_10209) );
ao12f01  g5400 ( .o(n10888), .a(n5658), .b(n6887), .c(x5548) );
oa12f01  g5401 ( .o(n3702), .a(n10888), .b(n6885_1), .c(n10887) );
in01f01  g5402 ( .o(n10890), .a(_net_10210) );
ao12f01  g5403 ( .o(n10891), .a(n5658), .b(n6887), .c(x5498) );
oa12f01  g5404 ( .o(n3707), .a(n10891), .b(n6885_1), .c(n10890) );
na03f01  g5405 ( .o(n10893), .a(n10045), .b(n6130), .c(_net_9385) );
no02f01  g5406 ( .o(n10894), .a(n6135), .b(n5658) );
na03f01  g5407 ( .o(n10895), .a(n10894), .b(n6140), .c(_net_9385) );
na03f01  g5408 ( .o(n10896), .a(n6136_1), .b(_net_9385), .c(x6599) );
no02f01  g5409 ( .o(n10897), .a(n6142), .b(n5658) );
oa12f01  g5410 ( .o(n10898), .a(n10897), .b(_net_9040), .c(_net_9385) );
na04f01  g5411 ( .o(n3712), .a(n10898), .b(n10896), .c(n10895), .d(n10893) );
in01f01  g5412 ( .o(n10900), .a(_net_131) );
oa12f01  g5413 ( .o(n3717), .a(n10900), .b(n9423), .c(n9419) );
no02f01  g5414 ( .o(n10902), .a(n9331), .b(_net_10372) );
na02f01  g5415 ( .o(n10903), .a(n9332), .b(n8183) );
oa12f01  g5416 ( .o(n10904), .a(n8200_1), .b(n9336), .c(_net_10372) );
ao12f01  g5417 ( .o(n10905), .a(n10904), .b(n9336), .c(_net_10372) );
ao12f01  g5418 ( .o(n10906), .a(n10905), .b(n8202), .c(_net_10372) );
oa12f01  g5419 ( .o(n3722), .a(n10906), .b(n10903), .c(n10902) );
ao12f01  g5420 ( .o(n10908), .a(n5658), .b(n7844), .c(net_249) );
ao22f01  g5421 ( .o(n10909), .a(n7847), .b(x4937), .c(n7846), .d(net_9811) );
na02f01  g5422 ( .o(n3727), .a(n10909), .b(n10908) );
na02f01  g5423 ( .o(n10911), .a(n6038), .b(_net_233) );
na02f01  g5424 ( .o(n10912), .a(n6037_1), .b(net_9862) );
ao22f01  g5425 ( .o(n10913), .a(n6044), .b(x5961), .c(n6042_1), .d(_net_10307) );
na04f01  g5426 ( .o(n3732), .a(n10913), .b(n10912), .c(n10911), .d(n6040) );
na02f01  g5427 ( .o(n10915), .a(n6020), .b(n6614_1) );
oa12f01  g5428 ( .o(n8762), .a(n10915), .b(n6020), .c(n7554) );
na02f01  g5429 ( .o(n10917), .a(n8762), .b(n7991) );
na02f01  g5430 ( .o(n10918), .a(n9463), .b(net_9523) );
ao12f01  g5431 ( .o(n10919), .a(n7999), .b(n10918), .c(n9620) );
in01f01  g5432 ( .o(n10920), .a(net_9523) );
oa12f01  g5433 ( .o(n10921), .a(x6599), .b(n8002), .c(n10920) );
no02f01  g5434 ( .o(n10922), .a(n10921), .b(n10919) );
na02f01  g5435 ( .o(n3737), .a(n10922), .b(n10917) );
in01f01  g5436 ( .o(n10924), .a(_net_9386) );
no02f01  g5437 ( .o(n10925), .a(n7446), .b(n10924) );
oa12f01  g5438 ( .o(n10926), .a(n10043), .b(n10925), .c(n10042) );
no02f01  g5439 ( .o(n10927), .a(_net_9040), .b(n10924) );
no03f01  g5440 ( .o(n10928), .a(n10924), .b(n6135), .c(n5658) );
ao22f01  g5441 ( .o(n10929), .a(n10928), .b(n6140), .c(n10927), .d(n10047) );
na02f01  g5442 ( .o(n3742), .a(n10929), .b(n10926) );
oa22f01  g5443 ( .o(n3750), .a(n7480_1), .b(n6785), .c(n7478), .d(n5573) );
ao22f01  g5444 ( .o(n10932), .a(n5842), .b(net_9671), .c(n5841), .d(net_109) );
na02f01  g5445 ( .o(n10933), .a(n5847), .b(net_9968) );
ao22f01  g5446 ( .o(n10934), .a(n5850), .b(net_9770), .c(n5849_1), .d(net_9869) );
na03f01  g5447 ( .o(n3763), .a(n10934), .b(n10933), .c(n10932) );
ao22f01  g5448 ( .o(n10936), .a(n5842), .b(net_9666), .c(n5841), .d(net_104) );
na02f01  g5449 ( .o(n10937), .a(n5847), .b(net_9963) );
ao22f01  g5450 ( .o(n10938), .a(n5850), .b(net_9765), .c(n5849_1), .d(net_9864) );
na03f01  g5451 ( .o(n3768), .a(n10938), .b(n10937), .c(n10936) );
no02f01  g5452 ( .o(n10940), .a(n9894), .b(_net_10229) );
na02f01  g5453 ( .o(n10941), .a(n10940), .b(n9220) );
in01f01  g5454 ( .o(n10942), .a(n10940) );
na02f01  g5455 ( .o(n10943), .a(n10942), .b(_net_10230) );
na02f01  g5456 ( .o(n3773), .a(n10943), .b(n10941) );
oa22f01  g5457 ( .o(n3778), .a(n5907), .b(n5833), .c(n5905), .d(n5612) );
na02f01  g5458 ( .o(n10946), .a(n5753_1), .b(_net_10120) );
na02f01  g5459 ( .o(n3787), .a(n10946), .b(n5755) );
in01f01  g5460 ( .o(n10948), .a(n6746) );
in01f01  g5461 ( .o(n10949), .a(_net_10149) );
in01f01  g5462 ( .o(n10950), .a(_net_10148) );
no02f01  g5463 ( .o(n10951), .a(n10950), .b(_net_9736) );
no02f01  g5464 ( .o(n10952), .a(_net_10148), .b(n8661) );
in01f01  g5465 ( .o(n10953), .a(n10952) );
no02f01  g5466 ( .o(n10954), .a(n10379), .b(_net_10147) );
ao12f01  g5467 ( .o(n10955), .a(n6737), .b(n6734), .c(n6719) );
in01f01  g5468 ( .o(n10956), .a(n10955) );
no02f01  g5469 ( .o(n10957), .a(n8532), .b(_net_10146) );
no02f01  g5470 ( .o(n10958), .a(n8525), .b(_net_10145) );
no03f01  g5471 ( .o(n10959), .a(n10958), .b(n10957), .c(n10956) );
in01f01  g5472 ( .o(n10960), .a(n10958) );
in01f01  g5473 ( .o(n10961), .a(_net_10145) );
no02f01  g5474 ( .o(n10962), .a(_net_9733), .b(n10961) );
ao12f01  g5475 ( .o(n10963), .a(n10962), .b(n10960), .c(n6739) );
no02f01  g5476 ( .o(n10964), .a(n10963), .b(n10957) );
in01f01  g5477 ( .o(n10965), .a(_net_10146) );
no02f01  g5478 ( .o(n10966), .a(_net_9734), .b(n10965) );
in01f01  g5479 ( .o(n10967), .a(_net_10147) );
no02f01  g5480 ( .o(n10968), .a(_net_9735), .b(n10967) );
no02f01  g5481 ( .o(n10969), .a(n10968), .b(n10966) );
ao12f01  g5482 ( .o(n10970), .a(n10969), .b(n10954), .c(_net_9735) );
no02f01  g5483 ( .o(n10971), .a(n10970), .b(n10964) );
in01f01  g5484 ( .o(n10972), .a(n10971) );
no02f01  g5485 ( .o(n10973), .a(n10972), .b(n10959) );
na02f01  g5486 ( .o(n10974), .a(n10970), .b(_net_10147) );
oa12f01  g5487 ( .o(n10975), .a(n10974), .b(n10973), .c(n10954) );
ao12f01  g5488 ( .o(n10976), .a(n10951), .b(n10975), .c(n10953) );
na02f01  g5489 ( .o(n10977), .a(n10976), .b(n10949) );
in01f01  g5490 ( .o(n10978), .a(n10977) );
no02f01  g5491 ( .o(n10979), .a(n10976), .b(n10949) );
oa12f01  g5492 ( .o(n10980), .a(n10948), .b(n10979), .c(n10978) );
no02f01  g5493 ( .o(n10981), .a(n10961), .b(n6738_1) );
in01f01  g5494 ( .o(n10982), .a(n10981) );
no02f01  g5495 ( .o(n10983), .a(n10982), .b(n6755) );
in01f01  g5496 ( .o(n10984), .a(n10983) );
no02f01  g5497 ( .o(n10985), .a(n10984), .b(n10965) );
in01f01  g5498 ( .o(n10986), .a(n10985) );
no02f01  g5499 ( .o(n10987), .a(n10986), .b(n10967) );
in01f01  g5500 ( .o(n10988), .a(n10987) );
no02f01  g5501 ( .o(n10989), .a(n10988), .b(n10950) );
in01f01  g5502 ( .o(n10990), .a(n10989) );
no02f01  g5503 ( .o(n10991), .a(n10990), .b(n10949) );
in01f01  g5504 ( .o(n10992), .a(n10991) );
ao12f01  g5505 ( .o(n10993), .a(n10398), .b(n10990), .c(n10949) );
ao22f01  g5506 ( .o(n10994), .a(n10993), .b(n10992), .c(n6760), .d(_net_10149) );
na02f01  g5507 ( .o(n3796), .a(n10994), .b(n10980) );
in01f01  g5508 ( .o(n10996), .a(x682) );
oa22f01  g5509 ( .o(n10997), .a(n10174), .b(net_9270), .c(n10158), .d(_net_9309) );
ao12f01  g5510 ( .o(n10998), .a(n10997), .b(n10171), .c(n7095_1) );
oa12f01  g5511 ( .o(n10999), .a(n10998), .b(n10170), .c(_net_9363) );
ao12f01  g5512 ( .o(n11000), .a(n10999), .b(n10163), .c(n7192_1) );
oa22f01  g5513 ( .o(n3801), .a(n11000), .b(n10157), .c(n10155), .d(n10996) );
na02f01  g5514 ( .o(n11002), .a(n6038), .b(_net_259) );
na02f01  g5515 ( .o(n11003), .a(n6037_1), .b(net_9888) );
ao22f01  g5516 ( .o(n11004), .a(n6044), .b(x4117), .c(n6042_1), .d(_net_10333) );
na04f01  g5517 ( .o(n3805), .a(n11004), .b(n11003), .c(n11002), .d(n6040) );
in01f01  g5518 ( .o(n11006), .a(net_10390) );
oa22f01  g5519 ( .o(n3810), .a(n10211), .b(n5615), .c(n10210), .d(n11006) );
na04f01  g5520 ( .o(n11008), .a(net_9221), .b(n9909), .c(n10509), .d(n9906) );
na04f01  g5521 ( .o(n11009), .a(net_9223), .b(net_9226), .c(n9908), .d(n9918) );
no02f01  g5522 ( .o(n3815), .a(n11009), .b(n11008) );
oa12f01  g5523 ( .o(n11011), .a(n7064), .b(n7001), .c(_net_10372) );
oa12f01  g5524 ( .o(n11012), .a(n11011), .b(n7002), .c(n7062) );
oa12f01  g5525 ( .o(n11013), .a(n11012), .b(n7063_1), .c(n7060) );
no02f01  g5526 ( .o(n11014), .a(n8931), .b(n9321) );
no02f01  g5527 ( .o(n11015), .a(_net_10335), .b(_net_10373) );
no02f01  g5528 ( .o(n11016), .a(n11015), .b(n11014) );
na02f01  g5529 ( .o(n11017), .a(n11016), .b(n11013) );
in01f01  g5530 ( .o(n11018), .a(n11013) );
in01f01  g5531 ( .o(n11019), .a(n11016) );
na02f01  g5532 ( .o(n11020), .a(n11019), .b(n11018) );
na02f01  g5533 ( .o(n3820), .a(n11020), .b(n11017) );
oa22f01  g5534 ( .o(n3825), .a(n5694), .b(n5719_1), .c(n5692), .d(n5649) );
oa22f01  g5535 ( .o(n3830), .a(n7738_1), .b(n7890), .c(n7736), .d(n9375) );
na02f01  g5536 ( .o(n11024), .a(n7358), .b(net_260) );
na02f01  g5537 ( .o(n11025), .a(n7352), .b(net_9691) );
ao22f01  g5538 ( .o(n11026), .a(n7357), .b(_net_10124), .c(n7353), .d(x4041) );
na04f01  g5539 ( .o(n3839), .a(n11026), .b(n11025), .c(n11024), .d(n7355_1) );
in01f01  g5540 ( .o(n3844), .a(n8108) );
na02f01  g5541 ( .o(n11029), .a(n6038), .b(net_250) );
na02f01  g5542 ( .o(n11030), .a(n6037_1), .b(net_9879) );
ao22f01  g5543 ( .o(n11031), .a(n6044), .b(x4851), .c(n6042_1), .d(_net_10324) );
na04f01  g5544 ( .o(n3849), .a(n11031), .b(n11030), .c(n11029), .d(n6040) );
ao12f01  g5545 ( .o(n11033), .a(n5658), .b(n5774), .c(x4520) );
oa12f01  g5546 ( .o(n3854), .a(n11033), .b(n5770), .c(n7044_1) );
na02f01  g5547 ( .o(n11035), .a(n6349), .b(n6326_1) );
oa22f01  g5548 ( .o(n3859), .a(n11035), .b(n6348), .c(n6349), .d(n8911) );
ao12f01  g5549 ( .o(n11037), .a(n5658), .b(n6532), .c(net_241) );
ao22f01  g5550 ( .o(n11038), .a(n6535), .b(x5498), .c(n6534), .d(net_10001) );
na02f01  g5551 ( .o(n3864), .a(n11038), .b(n11037) );
na02f01  g5552 ( .o(n11040), .a(n6349), .b(n6315) );
oa22f01  g5553 ( .o(n3869), .a(n11040), .b(n6348), .c(n6349), .d(n8896) );
in01f01  g5554 ( .o(n11042), .a(net_9230) );
no02f01  g5555 ( .o(n11043), .a(n7704_1), .b(n11042) );
no02f01  g5556 ( .o(n11044), .a(n7705), .b(net_9230) );
no03f01  g5557 ( .o(n3874), .a(n11044), .b(n11043), .c(n7703) );
in01f01  g5558 ( .o(n11046), .a(_net_10410) );
ao12f01  g5559 ( .o(n11047), .a(n5658), .b(n6052_1), .c(x6102) );
oa12f01  g5560 ( .o(n3879), .a(n11047), .b(n6048), .c(n11046) );
ao12f01  g5561 ( .o(n11049), .a(n5658), .b(n5678), .c(_net_234) );
ao22f01  g5562 ( .o(n11050), .a(n5681_1), .b(x5901), .c(n5680), .d(net_9697) );
na02f01  g5563 ( .o(n3884), .a(n11050), .b(n11049) );
ao12f01  g5564 ( .o(n11052), .a(n5658), .b(n5678), .c(net_237) );
ao22f01  g5565 ( .o(n11053), .a(n5681_1), .b(x5722), .c(n5680), .d(net_9700) );
na02f01  g5566 ( .o(n3889), .a(n11053), .b(n11052) );
no03f01  g5567 ( .o(n11055), .a(n7328), .b(n7322), .c(n7095_1) );
ao12f01  g5568 ( .o(n11056), .a(_net_9371), .b(n7332), .c(n7331_1) );
oa12f01  g5569 ( .o(n11057), .a(n10245), .b(n11056), .c(n11055) );
na03f01  g5570 ( .o(n11058), .a(n7332), .b(n7331_1), .c(_net_9371) );
oa12f01  g5571 ( .o(n11059), .a(n7095_1), .b(n7328), .c(n7322) );
na03f01  g5572 ( .o(n11060), .a(n11059), .b(n11058), .c(n10248) );
ao12f01  g5573 ( .o(n11061), .a(n10260), .b(n11060), .c(n11057) );
ao12f01  g5574 ( .o(n11062), .a(n10248), .b(n11059), .c(n11058) );
no03f01  g5575 ( .o(n11063), .a(n11056), .b(n11055), .c(n10245) );
no03f01  g5576 ( .o(n11064), .a(n11063), .b(n11062), .c(n10259) );
oa12f01  g5577 ( .o(n11065), .a(n6148), .b(n11064), .c(n11061) );
ao12f01  g5578 ( .o(n11066), .a(n6131_1), .b(n6147), .c(_net_9363) );
na02f01  g5579 ( .o(n3894), .a(n11066), .b(n11065) );
ao22f01  g5580 ( .o(n11068), .a(n5842), .b(net_9754), .c(n5841), .d(_net_190) );
na02f01  g5581 ( .o(n11069), .a(n5847), .b(net_10051) );
ao22f01  g5582 ( .o(n11070), .a(n5850), .b(net_9853), .c(n5849_1), .d(net_9952) );
na03f01  g5583 ( .o(n3899), .a(n11070), .b(n11069), .c(n11068) );
in01f01  g5584 ( .o(n11072), .a(net_9747) );
no02f01  g5585 ( .o(n11073), .a(n6976_1), .b(n5658) );
oa12f01  g5586 ( .o(n11074), .a(n11073), .b(n7366), .c(x4587) );
oa12f01  g5587 ( .o(n3904), .a(n11074), .b(n6977), .c(n11072) );
oa22f01  g5588 ( .o(n3909), .a(n7480_1), .b(n6595), .c(n7478), .d(n5576) );
in01f01  g5589 ( .o(n11077), .a(n8961) );
na03f01  g5590 ( .o(n11078), .a(n8965), .b(n8962), .c(n11077) );
oa12f01  g5591 ( .o(n11079), .a(n8963), .b(n8964), .c(n8961) );
na02f01  g5592 ( .o(n3914), .a(n11079), .b(n11078) );
na02f01  g5593 ( .o(n11081), .a(net_114), .b(_net_9606) );
ao12f01  g5594 ( .o(n11082), .a(n7543_1), .b(n7624), .c(n7512) );
no02f01  g5595 ( .o(n11083), .a(n11082), .b(net_9559) );
no02f01  g5596 ( .o(n11084), .a(n7636_1), .b(n7626_1) );
no03f01  g5597 ( .o(n11085), .a(n11084), .b(n7543_1), .c(n7625) );
oa12f01  g5598 ( .o(n11086), .a(n7500), .b(n11085), .c(n11083) );
na02f01  g5599 ( .o(n3923), .a(n11086), .b(n11081) );
no02f01  g5600 ( .o(n11088), .a(n7871_1), .b(_net_10458) );
no02f01  g5601 ( .o(n11089), .a(n9705), .b(n11088) );
oa12f01  g5602 ( .o(n11090), .a(n11089), .b(n9713), .c(n9704) );
no03f01  g5603 ( .o(n11091), .a(n11089), .b(n9713), .c(n9704) );
no02f01  g5604 ( .o(n11092), .a(n11091), .b(n7875) );
na02f01  g5605 ( .o(n11093), .a(n11092), .b(n11090) );
no02f01  g5606 ( .o(n11094), .a(n9728), .b(_net_10458) );
no02f01  g5607 ( .o(n11095), .a(n11094), .b(n9730) );
ao22f01  g5608 ( .o(n11096), .a(n11095), .b(n7450), .c(n7453), .d(_net_10458) );
na02f01  g5609 ( .o(n3928), .a(n11096), .b(n11093) );
in01f01  g5610 ( .o(n11098), .a(x3645) );
no02f01  g5611 ( .o(n3942), .a(n11098), .b(n5658) );
ao22f01  g5612 ( .o(n11100), .a(n5842), .b(net_9697), .c(n5841), .d(net_137) );
na02f01  g5613 ( .o(n11101), .a(n5847), .b(net_9994) );
ao22f01  g5614 ( .o(n11102), .a(n5850), .b(net_9796), .c(n5849_1), .d(net_9895) );
na03f01  g5615 ( .o(n3947), .a(n11102), .b(n11101), .c(n11100) );
in01f01  g5616 ( .o(n11104), .a(net_10498) );
oa22f01  g5617 ( .o(n3952), .a(n7467), .b(n5591), .c(n7465_1), .d(n11104) );
ao22f01  g5618 ( .o(n11106), .a(n6590), .b(net_10023), .c(n6580), .d(net_9793) );
ao22f01  g5619 ( .o(n11107), .a(n6584_1), .b(net_9761), .c(n6582), .d(net_9892) );
in01f01  g5620 ( .o(n11108), .a(n8051_1) );
ao22f01  g5621 ( .o(n11109), .a(n8047), .b(net_10059), .c(n8045), .d(net_224) );
oa12f01  g5622 ( .o(n11110), .a(n11109), .b(n11108), .c(n5520) );
na02f01  g5623 ( .o(n11111), .a(n8042), .b(net_10520) );
ao22f01  g5624 ( .o(n11112), .a(n6564), .b(net_10072), .c(n6562), .d(net_197) );
na02f01  g5625 ( .o(n11113), .a(n11112), .b(n11111) );
no02f01  g5626 ( .o(n11114), .a(n11113), .b(n11110) );
ao22f01  g5627 ( .o(n11115), .a(n6585), .b(net_9694), .c(n6573), .d(net_9860) );
ao22f01  g5628 ( .o(n11116), .a(n6605), .b(net_10294), .c(n6592), .d(net_10189) );
na02f01  g5629 ( .o(n11117), .a(n11116), .b(n11115) );
ao22f01  g5630 ( .o(n11118), .a(n6602), .b(net_9991), .c(n6572), .d(net_10399) );
ao22f01  g5631 ( .o(n11119), .a(n6603), .b(net_10504), .c(n6577), .d(net_9662) );
ao22f01  g5632 ( .o(n11120), .a(n6606), .b(net_9924), .c(n6597), .d(net_9726) );
ao22f01  g5633 ( .o(n11121), .a(n6599_1), .b(net_9825), .c(n6555), .d(net_9959) );
na04f01  g5634 ( .o(n11122), .a(n11121), .b(n11120), .c(n11119), .d(n11118) );
no02f01  g5635 ( .o(n11123), .a(n11122), .b(n11117) );
na04f01  g5636 ( .o(n3962), .a(n11123), .b(n11114), .c(n11107), .d(n11106) );
na02f01  g5637 ( .o(n11125), .a(n8017), .b(_net_9177) );
na02f01  g5638 ( .o(n11126), .a(_net_9178), .b(n1521) );
na02f01  g5639 ( .o(n3967), .a(n11126), .b(n11125) );
ao12f01  g5640 ( .o(n11128), .a(n5658), .b(n6160_1), .c(x4851) );
oa12f01  g5641 ( .o(n3972), .a(n11128), .b(n6159), .c(n3146) );
ao12f01  g5642 ( .o(n11130), .a(n7884), .b(n9756), .c(n7732) );
oa12f01  g5643 ( .o(n11131), .a(n7921_1), .b(n11130), .c(n7908) );
no02f01  g5644 ( .o(n11132), .a(n7884), .b(n7732) );
oa12f01  g5645 ( .o(n11133), .a(_net_9356), .b(n8754), .c(net_9151) );
no02f01  g5646 ( .o(n11134), .a(n7734_1), .b(n7884) );
ao22f01  g5647 ( .o(n11135), .a(n11134), .b(n9772), .c(n9774), .d(_net_9356) );
oa12f01  g5648 ( .o(n11136), .a(n11135), .b(n11133), .c(n9769) );
ao12f01  g5649 ( .o(n11137), .a(n11136), .b(n11132), .c(n9766) );
oa12f01  g5650 ( .o(n3980), .a(n11137), .b(n11131), .c(n9760) );
na02f01  g5651 ( .o(n11139), .a(n6056), .b(net_245) );
na02f01  g5652 ( .o(n11140), .a(n6055), .b(net_9973) );
ao22f01  g5653 ( .o(n11141), .a(n6062_1), .b(x5225), .c(n6060), .d(_net_10424) );
na04f01  g5654 ( .o(n3985), .a(n11141), .b(n11140), .c(n11139), .d(n6058) );
in01f01  g5655 ( .o(n11143), .a(_net_9352) );
no02f01  g5656 ( .o(n3990), .a(n8637), .b(n11143) );
in01f01  g5657 ( .o(n11145), .a(_net_9643) );
no03f01  g5658 ( .o(n11146), .a(n9540), .b(n7966), .c(n11145) );
na03f01  g5659 ( .o(n11147), .a(n9542), .b(_net_9643), .c(_net_9641) );
na02f01  g5660 ( .o(n11148), .a(n9495), .b(_net_9643) );
no02f01  g5661 ( .o(n11149), .a(n9546), .b(n11145) );
oa22f01  g5662 ( .o(n11150), .a(n9791), .b(n11145), .c(_net_9250), .d(n9786) );
ao12f01  g5663 ( .o(n11151), .a(n11150), .b(n11149), .c(n8774) );
na03f01  g5664 ( .o(n11152), .a(n11151), .b(n11148), .c(n11147) );
oa12f01  g5665 ( .o(n11153), .a(x6599), .b(n11152), .c(n11146) );
no02f01  g5666 ( .o(n3994), .a(n11153), .b(n2827) );
in01f01  g5667 ( .o(n11155), .a(_net_10151) );
no03f01  g5668 ( .o(n11156), .a(n10977), .b(_net_10150), .c(n11155) );
no02f01  g5669 ( .o(n11157), .a(n10977), .b(_net_10150) );
oa12f01  g5670 ( .o(n11158), .a(n10948), .b(n11157), .c(_net_10151) );
na02f01  g5671 ( .o(n11159), .a(n10991), .b(_net_10150) );
in01f01  g5672 ( .o(n11160), .a(n11159) );
na02f01  g5673 ( .o(n11161), .a(n11160), .b(_net_10151) );
ao12f01  g5674 ( .o(n11162), .a(n10398), .b(n11159), .c(n11155) );
ao22f01  g5675 ( .o(n11163), .a(n11162), .b(n11161), .c(n6760), .d(_net_10151) );
oa12f01  g5676 ( .o(n3999), .a(n11163), .b(n11158), .c(n11156) );
na02f01  g5677 ( .o(n11165), .a(net_10186), .b(net_10194) );
ao22f01  g5678 ( .o(n11166), .a(net_10187), .b(net_10195), .c(net_10185), .d(net_10193) );
ao22f01  g5679 ( .o(n11167), .a(net_10182), .b(net_10189), .c(net_10185), .d(net_10192) );
ao22f01  g5680 ( .o(n11168), .a(net_10184), .b(net_10191), .c(net_10183), .d(net_10190) );
na04f01  g5681 ( .o(n4004), .a(n11168), .b(n11167), .c(n11166), .d(n11165) );
na02f01  g5682 ( .o(n11170), .a(n5755), .b(_net_10121) );
na02f01  g5683 ( .o(n4009), .a(n11170), .b(n5757) );
no02f01  g5684 ( .o(n11172), .a(n6713_1), .b(_net_9731) );
no02f01  g5685 ( .o(n11173), .a(n11172), .b(n6721) );
oa12f01  g5686 ( .o(n11174), .a(n11173), .b(n6733_1), .c(n6715) );
no03f01  g5687 ( .o(n11175), .a(n11173), .b(n6733_1), .c(n6715) );
no02f01  g5688 ( .o(n11176), .a(n11175), .b(n6746) );
na02f01  g5689 ( .o(n11177), .a(n11176), .b(n11174) );
no02f01  g5690 ( .o(n11178), .a(n6754), .b(_net_10143) );
no02f01  g5691 ( .o(n11179), .a(n11178), .b(n6756) );
ao22f01  g5692 ( .o(n11180), .a(n11179), .b(n6750), .c(n6760), .d(_net_10143) );
na02f01  g5693 ( .o(n4014), .a(n11180), .b(n11177) );
ao12f01  g5694 ( .o(n11182), .a(n5658), .b(n6875_1), .c(net_245) );
ao22f01  g5695 ( .o(n11183), .a(n6878), .b(x5225), .c(n6877), .d(net_9906) );
na02f01  g5696 ( .o(n4019), .a(n11183), .b(n11182) );
in01f01  g5697 ( .o(n11185), .a(_net_10109) );
ao12f01  g5698 ( .o(n11186), .a(n5658), .b(n6160_1), .c(x5225) );
oa12f01  g5699 ( .o(n4024), .a(n11186), .b(n6159), .c(n11185) );
in01f01  g5700 ( .o(n11188), .a(_net_10426) );
ao12f01  g5701 ( .o(n11189), .a(n5658), .b(n6052_1), .c(x5077) );
oa12f01  g5702 ( .o(n4029), .a(n11189), .b(n6048), .c(n11188) );
na02f01  g5703 ( .o(n11191), .a(_net_9296), .b(_net_9606) );
oa12f01  g5704 ( .o(n4034), .a(n11191), .b(_net_9606), .c(n9869) );
ao12f01  g5705 ( .o(n11193), .a(n5658), .b(n7844), .c(net_251) );
ao22f01  g5706 ( .o(n11194), .a(n7847), .b(x4781), .c(n7846), .d(net_9813) );
na02f01  g5707 ( .o(n4039), .a(n11194), .b(n11193) );
na02f01  g5708 ( .o(n11196), .a(n6038), .b(net_244) );
na02f01  g5709 ( .o(n11197), .a(n6037_1), .b(net_9873) );
ao22f01  g5710 ( .o(n11198), .a(n6044), .b(x5289), .c(n6042_1), .d(_net_10318) );
na04f01  g5711 ( .o(n4044), .a(n11198), .b(n11197), .c(n11196), .d(n6040) );
ao12f01  g5712 ( .o(n11200), .a(n5658), .b(n5774), .c(x4041) );
oa12f01  g5713 ( .o(n4049), .a(n11200), .b(n5770), .c(n7064) );
no02f01  g5714 ( .o(n11202), .a(n6808), .b(n6779) );
ao12f01  g5715 ( .o(n11203), .a(n6933), .b(n11202), .c(n6795) );
oa12f01  g5716 ( .o(n11204), .a(n11203), .b(n11202), .c(n6795) );
no02f01  g5717 ( .o(n11205), .a(n6834), .b(_net_10249) );
no02f01  g5718 ( .o(n11206), .a(n6835), .b(n6807) );
no02f01  g5719 ( .o(n11207), .a(n11206), .b(n11205) );
ao22f01  g5720 ( .o(n11208), .a(n11207), .b(n6175), .c(n6168), .d(_net_10249) );
na02f01  g5721 ( .o(n4054), .a(n11208), .b(n11204) );
in01f01  g5722 ( .o(n11210), .a(net_223) );
in01f01  g5723 ( .o(n11211), .a(net_222) );
no02f01  g5724 ( .o(n11212), .a(n10370), .b(n11211) );
in01f01  g5725 ( .o(n11213), .a(n11212) );
na02f01  g5726 ( .o(n11214), .a(n11213), .b(n11210) );
na02f01  g5727 ( .o(n11215), .a(n11212), .b(net_223) );
na02f01  g5728 ( .o(n11216), .a(n11215), .b(n11214) );
oa22f01  g5729 ( .o(n4059), .a(n11216), .b(n10367), .c(n10373), .d(n11210) );
na02f01  g5730 ( .o(n11218), .a(_net_178), .b(net_313) );
in01f01  g5731 ( .o(n11219), .a(n11218) );
no02f01  g5732 ( .o(n11220), .a(n5918), .b(n9549) );
in01f01  g5733 ( .o(n11221), .a(n11220) );
na02f01  g5734 ( .o(n11222), .a(_net_179), .b(net_313) );
in01f01  g5735 ( .o(n11223), .a(n11222) );
no03f01  g5736 ( .o(n11224), .a(n11223), .b(n11221), .c(n11219) );
no02f01  g5737 ( .o(n11225), .a(n11224), .b(n5921_1) );
in01f01  g5738 ( .o(n11226), .a(n11224) );
no02f01  g5739 ( .o(n11227), .a(n11226), .b(n5931_1) );
no02f01  g5740 ( .o(n11228), .a(n11227), .b(n11225) );
na02f01  g5741 ( .o(n11229), .a(n11224), .b(n5931_1) );
ao12f01  g5742 ( .o(n11230), .a(n7898_1), .b(n7904), .c(n7894) );
in01f01  g5743 ( .o(n11231), .a(_net_190) );
na02f01  g5744 ( .o(n11232), .a(n11223), .b(n11231) );
no02f01  g5745 ( .o(n11233), .a(n11232), .b(n11218) );
no03f01  g5746 ( .o(n11234), .a(n9551), .b(_net_188), .c(_net_189) );
in01f01  g5747 ( .o(n11235), .a(n11233) );
oa12f01  g5748 ( .o(n11236), .a(n11235), .b(n11222), .c(_net_189) );
no02f01  g5749 ( .o(n11237), .a(n9551), .b(_net_187) );
ao22f01  g5750 ( .o(n11238), .a(n11237), .b(n11236), .c(n11234), .d(n11233) );
oa22f01  g5751 ( .o(n4064), .a(n11238), .b(n11228), .c(n11230), .d(n11229) );
in01f01  g5752 ( .o(n11240), .a(_net_10441) );
ao12f01  g5753 ( .o(n11241), .a(n5658), .b(n6052_1), .c(x3889) );
oa12f01  g5754 ( .o(n4069), .a(n11241), .b(n6048), .c(n11240) );
in01f01  g5755 ( .o(n11243), .a(net_10404) );
in01f01  g5756 ( .o(n11244), .a(net_10398) );
na02f01  g5757 ( .o(n11245), .a(n11244), .b(x6599) );
na02f01  g5758 ( .o(n11246), .a(net_263), .b(net_10385) );
ao12f01  g5759 ( .o(n4074), .a(n11245), .b(n11246), .c(n11243) );
ao12f01  g5760 ( .o(n11248), .a(n5658), .b(n7844), .c(net_245) );
ao22f01  g5761 ( .o(n11249), .a(n7847), .b(x5225), .c(n7846), .d(net_9807) );
na02f01  g5762 ( .o(n4079), .a(n11249), .b(n11248) );
in01f01  g5763 ( .o(n11251), .a(_net_10316) );
ao12f01  g5764 ( .o(n11252), .a(n5658), .b(n5774), .c(x5427) );
oa12f01  g5765 ( .o(n4093), .a(n11252), .b(n5770), .c(n11251) );
ao12f01  g5766 ( .o(n11254), .a(n7546), .b(n6028_1), .c(n6634_1) );
oa12f01  g5767 ( .o(n4098), .a(n11254), .b(n6022), .c(n8466) );
in01f01  g5768 ( .o(n11256), .a(net_9852) );
oa12f01  g5769 ( .o(n11257), .a(x6599), .b(n8828), .c(n7841) );
na02f01  g5770 ( .o(n11258), .a(n8830), .b(net_10280) );
oa22f01  g5771 ( .o(n4103), .a(n11258), .b(n8827), .c(n11257), .d(n11256) );
na04f01  g5772 ( .o(n11260), .a(n8784), .b(n8753), .c(n9786), .d(_net_9637) );
no04f01  g5773 ( .o(n11261), .a(n11260), .b(n10494), .c(_net_9640), .d(_net_9639) );
ao12f01  g5774 ( .o(n11262), .a(net_9571), .b(_net_9573), .c(net_9647) );
oa12f01  g5775 ( .o(n4112), .a(n11262), .b(n11261), .c(n8743) );
oa22f01  g5776 ( .o(n4124), .a(n7367), .b(n6958_1), .c(n7365_1), .d(n5600) );
no02f01  g5777 ( .o(n11265), .a(n8225), .b(n8220) );
in01f01  g5778 ( .o(n11266), .a(n11265) );
na02f01  g5779 ( .o(n11267), .a(n11266), .b(n8233) );
na02f01  g5780 ( .o(n11268), .a(n11265), .b(n8232) );
na02f01  g5781 ( .o(n4129), .a(n11268), .b(n11267) );
ao12f01  g5782 ( .o(n11270), .a(n5658), .b(n5678), .c(_net_255) );
ao22f01  g5783 ( .o(n11271), .a(n5681_1), .b(x4449), .c(n5680), .d(net_9718) );
na02f01  g5784 ( .o(n4137), .a(n11271), .b(n11270) );
ao22f01  g5785 ( .o(n11273), .a(n5702), .b(x2477), .c(n5701), .d(_net_9402) );
oa12f01  g5786 ( .o(n4142), .a(n11273), .b(n5700_1), .c(n8114) );
in01f01  g5787 ( .o(n11275), .a(net_10297) );
na02f01  g5788 ( .o(n11276), .a(n9799), .b(net_10280) );
ao12f01  g5789 ( .o(n4147), .a(n5911), .b(n11276), .c(n11275) );
ao12f01  g5790 ( .o(n11278), .a(n5658), .b(n6875_1), .c(net_242) );
ao22f01  g5791 ( .o(n11279), .a(n6878), .b(x5427), .c(n6877), .d(net_9903) );
na02f01  g5792 ( .o(n4156), .a(n11279), .b(n11278) );
ao22f01  g5793 ( .o(n11281), .a(n5842), .b(net_9676), .c(n5841), .d(net_114) );
na02f01  g5794 ( .o(n11282), .a(n5847), .b(net_9973) );
ao22f01  g5795 ( .o(n11283), .a(n5850), .b(net_9775), .c(n5849_1), .d(net_9874) );
na03f01  g5796 ( .o(n4161), .a(n11283), .b(n11282), .c(n11281) );
oa22f01  g5797 ( .o(n4165), .a(n7480_1), .b(n6801_1), .c(n7478), .d(n5618) );
no02f01  g5798 ( .o(n11286), .a(n6806_1), .b(n6802) );
no03f01  g5799 ( .o(n11287), .a(n11286), .b(n6808), .c(n6797) );
oa12f01  g5800 ( .o(n11288), .a(n11286), .b(n6808), .c(n6797) );
na02f01  g5801 ( .o(n11289), .a(n11288), .b(n6177_1) );
oa12f01  g5802 ( .o(n11290), .a(n6175), .b(n11206), .c(_net_10250) );
ao12f01  g5803 ( .o(n11291), .a(n11290), .b(n11206), .c(_net_10250) );
ao12f01  g5804 ( .o(n11292), .a(n11291), .b(n6168), .c(_net_10250) );
oa12f01  g5805 ( .o(n4170), .a(n11292), .b(n11289), .c(n11287) );
in01f01  g5806 ( .o(n11294), .a(net_9841) );
oa22f01  g5807 ( .o(n4175), .a(n7480_1), .b(n11294), .c(n7478), .d(n5591) );
ao22f01  g5808 ( .o(n11296), .a(n5842), .b(net_9683), .c(n5841), .d(_net_121) );
na02f01  g5809 ( .o(n11297), .a(n5847), .b(net_9980) );
ao22f01  g5810 ( .o(n11298), .a(n5850), .b(net_9782), .c(n5849_1), .d(net_9881) );
na03f01  g5811 ( .o(n4180), .a(n11298), .b(n11297), .c(n11296) );
in01f01  g5812 ( .o(n11300), .a(net_10093) );
na02f01  g5813 ( .o(n11301), .a(_net_10094), .b(n11300) );
ao12f01  g5814 ( .o(n4185), .a(n6155_1), .b(n11301), .c(n10701) );
na02f01  g5815 ( .o(n11303), .a(n7398_1), .b(_net_10429) );
na02f01  g5816 ( .o(n4190), .a(n11303), .b(n8326) );
oa22f01  g5817 ( .o(n11305), .a(n6727), .b(_net_8846), .c(_net_10164), .d(n6729) );
na02f01  g5818 ( .o(n11306), .a(_net_10164), .b(n6729) );
oa22f01  g5819 ( .o(n11307), .a(n6723_1), .b(_net_10165), .c(_net_10166), .d(n6720) );
ao12f01  g5820 ( .o(n11308), .a(n11307), .b(n11306), .c(n11305) );
in01f01  g5821 ( .o(n11309), .a(_net_10166) );
oa12f01  g5822 ( .o(n11310), .a(_net_10165), .b(_net_10166), .c(n6720) );
oa22f01  g5823 ( .o(n11311), .a(n11310), .b(_net_9730), .c(n11309), .d(_net_9731) );
no02f01  g5824 ( .o(n11312), .a(n11311), .b(n11308) );
oa22f01  g5825 ( .o(n11313), .a(n10379), .b(net_10170), .c(net_10169), .d(n8532) );
oa22f01  g5826 ( .o(n11314), .a(_net_10167), .b(n6736), .c(n8525), .d(_net_10168) );
no03f01  g5827 ( .o(n11315), .a(n11314), .b(n11313), .c(n11312) );
in01f01  g5828 ( .o(n11316), .a(_net_10168) );
in01f01  g5829 ( .o(n11317), .a(_net_10167) );
ao12f01  g5830 ( .o(n11318), .a(n11317), .b(_net_9733), .c(n11316) );
ao22f01  g5831 ( .o(n11319), .a(n11318), .b(n6736), .c(n8525), .d(_net_10168) );
oa12f01  g5832 ( .o(n11320), .a(net_10169), .b(n10379), .c(net_10170) );
no02f01  g5833 ( .o(n11321), .a(n11320), .b(_net_9734) );
ao12f01  g5834 ( .o(n11322), .a(n11321), .b(n10379), .c(net_10170) );
oa12f01  g5835 ( .o(n11323), .a(n11322), .b(n11319), .c(n11313) );
oa22f01  g5836 ( .o(n11324), .a(n11323), .b(n11315), .c(_net_10171), .d(n8661) );
na02f01  g5837 ( .o(n11325), .a(_net_10171), .b(n8661) );
no03f01  g5838 ( .o(n11326), .a(_net_8819), .b(net_8818), .c(net_8838) );
na03f01  g5839 ( .o(n4195), .a(n11326), .b(n11325), .c(n11324) );
na02f01  g5840 ( .o(n11328), .a(n8947), .b(_net_10334) );
na02f01  g5841 ( .o(n4200), .a(n11328), .b(n8950) );
in01f01  g5842 ( .o(n11330), .a(n10314) );
no02f01  g5843 ( .o(n11331), .a(n10313), .b(n9048) );
oa12f01  g5844 ( .o(n11332), .a(n7431), .b(n11331), .c(n11330) );
no02f01  g5845 ( .o(n11333), .a(n9733), .b(n9037) );
in01f01  g5846 ( .o(n11334), .a(n11333) );
no02f01  g5847 ( .o(n11335), .a(n11334), .b(n10298) );
in01f01  g5848 ( .o(n11336), .a(n11335) );
no02f01  g5849 ( .o(n11337), .a(n11336), .b(n9048) );
in01f01  g5850 ( .o(n11338), .a(n11337) );
ao12f01  g5851 ( .o(n11339), .a(n7451_1), .b(n11336), .c(n9048) );
ao22f01  g5852 ( .o(n11340), .a(n11339), .b(n11338), .c(n7453), .d(_net_10464) );
na02f01  g5853 ( .o(n4205), .a(n11340), .b(n11332) );
in01f01  g5854 ( .o(n11342), .a(net_9228) );
in01f01  g5855 ( .o(n11343), .a(net_9231) );
no04f01  g5856 ( .o(n4210), .a(n11343), .b(n11042), .c(n11342), .d(net_9229) );
ao12f01  g5857 ( .o(n11345), .a(n8579), .b(n5922), .c(net_9568) );
in01f01  g5858 ( .o(n11346), .a(n11345) );
no02f01  g5859 ( .o(n4220), .a(n11346), .b(n5935_1) );
ao22f01  g5860 ( .o(n11348), .a(n5842), .b(net_9721), .c(n5841), .d(_net_161) );
na02f01  g5861 ( .o(n11349), .a(n5847), .b(net_10018) );
ao22f01  g5862 ( .o(n11350), .a(n5850), .b(net_9820), .c(n5849_1), .d(net_9919) );
na03f01  g5863 ( .o(n4225), .a(n11350), .b(n11349), .c(n11348) );
in01f01  g5864 ( .o(n11352), .a(net_10183) );
oa22f01  g5865 ( .o(n4230), .a(n7956), .b(n5591), .c(n7955), .d(n11352) );
oa12f01  g5866 ( .o(n11354), .a(n10963), .b(n10958), .c(n10956) );
no02f01  g5867 ( .o(n11355), .a(n10966), .b(n10957) );
ao12f01  g5868 ( .o(n11356), .a(n6746), .b(n11355), .c(n11354) );
oa12f01  g5869 ( .o(n11357), .a(n11356), .b(n11355), .c(n11354) );
na02f01  g5870 ( .o(n11358), .a(n10984), .b(n10965) );
no02f01  g5871 ( .o(n11359), .a(n10985), .b(n10398) );
ao22f01  g5872 ( .o(n11360), .a(n11359), .b(n11358), .c(n6760), .d(_net_10146) );
na02f01  g5873 ( .o(n4235), .a(n11360), .b(n11357) );
in01f01  g5874 ( .o(n11362), .a(net_9529) );
na02f01  g5875 ( .o(n11363), .a(n9468), .b(n11362) );
na02f01  g5876 ( .o(n11364), .a(n9469), .b(net_9529) );
ao12f01  g5877 ( .o(n11365), .a(n7999), .b(n11364), .c(n11363) );
oa12f01  g5878 ( .o(n11366), .a(x6599), .b(n8002), .c(n11362) );
no02f01  g5879 ( .o(n11367), .a(n11366), .b(n11365) );
oa12f01  g5880 ( .o(n4240), .a(n11367), .b(n10744), .c(n9454) );
ao12f01  g5881 ( .o(n11369), .a(n5658), .b(n6875_1), .c(_net_231) );
ao22f01  g5882 ( .o(n11370), .a(n6878), .b(x6102), .c(n6877), .d(net_9892) );
na02f01  g5883 ( .o(n4245), .a(n11370), .b(n11369) );
no02f01  g5884 ( .o(n11372), .a(_net_10534), .b(n5658) );
oa12f01  g5885 ( .o(n4250), .a(n11372), .b(n10629), .c(n5495_1) );
no02f01  g5886 ( .o(n11374), .a(n10472), .b(n10347) );
no02f01  g5887 ( .o(n11375), .a(n10471), .b(n10344) );
no02f01  g5888 ( .o(n11376), .a(net_9156), .b(net_9155) );
no02f01  g5889 ( .o(n11377), .a(n9168), .b(n7731) );
no02f01  g5890 ( .o(n11378), .a(n11377), .b(n11376) );
in01f01  g5891 ( .o(n11379), .a(n11378) );
no02f01  g5892 ( .o(n11380), .a(n11379), .b(net_9154) );
no02f01  g5893 ( .o(n11381), .a(n11378), .b(n8984) );
no04f01  g5894 ( .o(n11382), .a(n11381), .b(n11380), .c(n11375), .d(n11374) );
no02f01  g5895 ( .o(n11383), .a(n11375), .b(n11374) );
no02f01  g5896 ( .o(n11384), .a(n11381), .b(n11380) );
no02f01  g5897 ( .o(n11385), .a(n11384), .b(n11383) );
no02f01  g5898 ( .o(n11386), .a(n11385), .b(n11382) );
in01f01  g5899 ( .o(n11387), .a(n11386) );
no02f01  g5900 ( .o(n11388), .a(n11387), .b(_net_9320) );
no02f01  g5901 ( .o(n11389), .a(n11386), .b(n8332) );
no02f01  g5902 ( .o(n11390), .a(_net_9321), .b(_net_9322) );
no02f01  g5903 ( .o(n11391), .a(n8763), .b(n8658) );
no02f01  g5904 ( .o(n11392), .a(n11391), .b(n11390) );
in01f01  g5905 ( .o(n11393), .a(n11392) );
no03f01  g5906 ( .o(n11394), .a(n11393), .b(n11389), .c(n11388) );
no02f01  g5907 ( .o(n11395), .a(n11389), .b(n11388) );
no02f01  g5908 ( .o(n11396), .a(n11392), .b(n11395) );
no02f01  g5909 ( .o(n11397), .a(n11396), .b(n11394) );
no02f01  g5910 ( .o(n11398), .a(n10477), .b(n8989) );
no02f01  g5911 ( .o(n11399), .a(n10468), .b(n8983) );
no02f01  g5912 ( .o(n11400), .a(n11399), .b(n11398) );
no02f01  g5913 ( .o(n11401), .a(n11400), .b(n11397) );
na02f01  g5914 ( .o(n11402), .a(n11400), .b(n11397) );
na02f01  g5915 ( .o(n11403), .a(n11402), .b(n8638) );
ao12f01  g5916 ( .o(n11404), .a(n7883), .b(n8637), .c(_net_9312) );
oa12f01  g5917 ( .o(n4259), .a(n11404), .b(n11403), .c(n11401) );
no02f01  g5918 ( .o(n11406), .a(n11235), .b(n11221) );
in01f01  g5919 ( .o(n11407), .a(n11406) );
no02f01  g5920 ( .o(n11408), .a(n11218), .b(n11231) );
in01f01  g5921 ( .o(n11409), .a(n11408) );
no03f01  g5922 ( .o(n11410), .a(n11409), .b(n11222), .c(n11221) );
no02f01  g5923 ( .o(n11411), .a(n11410), .b(n5921_1) );
in01f01  g5924 ( .o(n11412), .a(n11411) );
na03f01  g5925 ( .o(n11413), .a(n11223), .b(n11218), .c(_net_185) );
na03f01  g5926 ( .o(n11414), .a(n11223), .b(_net_189), .c(_net_185) );
ao12f01  g5927 ( .o(n11415), .a(n5918), .b(n11414), .c(n11413) );
no02f01  g5928 ( .o(n11416), .a(n11415), .b(n5921_1) );
no03f01  g5929 ( .o(n11417), .a(n11416), .b(n11412), .c(n11407) );
no02f01  g5930 ( .o(n11418), .a(n11416), .b(n11412) );
no02f01  g5931 ( .o(n11419), .a(n11411), .b(n11406) );
no02f01  g5932 ( .o(n11420), .a(n11412), .b(n11407) );
no03f01  g5933 ( .o(n11421), .a(n11420), .b(n11419), .c(n11418) );
in01f01  g5934 ( .o(n11422), .a(n11421) );
no03f01  g5935 ( .o(n11423), .a(n11416), .b(n11411), .c(n11406) );
in01f01  g5936 ( .o(n11424), .a(n11423) );
na03f01  g5937 ( .o(n11425), .a(n11424), .b(n11422), .c(n7902_1) );
in01f01  g5938 ( .o(n11426), .a(_net_189) );
in01f01  g5939 ( .o(n11427), .a(net_186) );
na04f01  g5940 ( .o(n11428), .a(n11223), .b(n11427), .c(n5918), .d(n11426) );
no03f01  g5941 ( .o(n11429), .a(_net_189), .b(_net_187), .c(_net_185) );
no03f01  g5942 ( .o(n11430), .a(_net_188), .b(_net_189), .c(_net_185) );
no02f01  g5943 ( .o(n11431), .a(n11430), .b(n11429) );
oa12f01  g5944 ( .o(n11432), .a(n11431), .b(n11428), .c(n11408) );
no02f01  g5945 ( .o(n11433), .a(n5926_1), .b(n11426) );
in01f01  g5946 ( .o(n11434), .a(n11433) );
no02f01  g5947 ( .o(n11435), .a(n11434), .b(net_9622) );
no02f01  g5948 ( .o(n11436), .a(n11435), .b(n11424) );
ao12f01  g5949 ( .o(n11437), .a(n11436), .b(n11432), .c(n11421) );
oa12f01  g5950 ( .o(n4264), .a(n11437), .b(n11425), .c(n11417) );
no02f01  g5951 ( .o(n11439), .a(n9080), .b(n9079) );
ao12f01  g5952 ( .o(n11440), .a(n8184), .b(n11439), .c(n9120) );
oa12f01  g5953 ( .o(n11441), .a(n11440), .b(n11439), .c(n9120) );
in01f01  g5954 ( .o(n11442), .a(n9141) );
no02f01  g5955 ( .o(n11443), .a(n9140), .b(_net_10358) );
no03f01  g5956 ( .o(n11444), .a(n11443), .b(n11442), .c(n9144) );
ao12f01  g5957 ( .o(n11445), .a(n11444), .b(n8202), .c(_net_10358) );
na02f01  g5958 ( .o(n4269), .a(n11445), .b(n11441) );
ao22f01  g5959 ( .o(n11447), .a(n5842), .b(net_9675), .c(n5841), .d(net_113) );
na02f01  g5960 ( .o(n11448), .a(n5847), .b(net_9972) );
ao22f01  g5961 ( .o(n11449), .a(n5850), .b(net_9774), .c(n5849_1), .d(net_9873) );
na03f01  g5962 ( .o(n4274), .a(n11449), .b(n11448), .c(n11447) );
no03f01  g5963 ( .o(n11451), .a(n11235), .b(net_186), .c(n11426) );
na02f01  g5964 ( .o(n11452), .a(n11232), .b(n11219) );
na02f01  g5965 ( .o(n11453), .a(n11452), .b(n11237) );
no04f01  g5966 ( .o(n11454), .a(n11413), .b(net_186), .c(_net_188), .d(_net_189) );
na02f01  g5967 ( .o(n11455), .a(_net_189), .b(n9549) );
ao12f01  g5968 ( .o(n11456), .a(n11455), .b(_net_188), .c(_net_187) );
no02f01  g5969 ( .o(n11457), .a(n11456), .b(n11454) );
na02f01  g5970 ( .o(n11458), .a(n11457), .b(n11453) );
ao12f01  g5971 ( .o(n11459), .a(n11458), .b(n11451), .c(n5918) );
na02f01  g5972 ( .o(n11460), .a(n5926_1), .b(_net_190) );
na02f01  g5973 ( .o(n11461), .a(n11460), .b(n11434) );
no03f01  g5974 ( .o(n11462), .a(n11224), .b(n5931_1), .c(net_9622) );
no03f01  g5975 ( .o(n11463), .a(n11229), .b(n7906_1), .c(n7899) );
ao12f01  g5976 ( .o(n11464), .a(n11463), .b(n11462), .c(n11461) );
oa12f01  g5977 ( .o(n4283), .a(n11464), .b(n11459), .c(n11228) );
oa12f01  g5978 ( .o(n11466), .a(n7732), .b(n10524), .c(net_9657) );
ao12f01  g5979 ( .o(n4288), .a(n11466), .b(n10524), .c(net_9657) );
no02f01  g5980 ( .o(n11468), .a(n6561_1), .b(n11211) );
ao22f01  g5981 ( .o(n11469), .a(n11468), .b(n6558), .c(n6585), .d(net_9724) );
ao22f01  g5982 ( .o(n11470), .a(n6599_1), .b(net_9854), .c(n6584_1), .d(net_9791) );
ao22f01  g5983 ( .o(n11471), .a(n6573), .b(net_9890), .c(n6555), .d(net_9989) );
na02f01  g5984 ( .o(n11472), .a(n6582), .b(net_9922) );
ao22f01  g5985 ( .o(n11473), .a(n6580), .b(net_9823), .c(n6577), .d(net_9692) );
na02f01  g5986 ( .o(n11474), .a(n11473), .b(n11472) );
in01f01  g5987 ( .o(n11475), .a(net_9755) );
in01f01  g5988 ( .o(n11476), .a(net_9953) );
oa22f01  g5989 ( .o(n11477), .a(n6966_1), .b(n11476), .c(n6598), .d(n11475) );
in01f01  g5990 ( .o(n11478), .a(net_10021) );
in01f01  g5991 ( .o(n11479), .a(net_10052) );
oa22f01  g5992 ( .o(n11480), .a(n6959), .b(n11478), .c(n6591), .d(n11479) );
no03f01  g5993 ( .o(n11481), .a(n11480), .b(n11477), .c(n11474) );
na04f01  g5994 ( .o(n4298), .a(n11481), .b(n11471), .c(n11470), .d(n11469) );
na02f01  g5995 ( .o(n11483), .a(n7937), .b(net_246) );
na02f01  g5996 ( .o(n11484), .a(n7936), .b(net_9776) );
ao22f01  g5997 ( .o(n11485), .a(n7943), .b(_net_10215), .c(n7942), .d(x5143) );
na04f01  g5998 ( .o(n4303), .a(n11485), .b(n11484), .c(n11483), .d(n7939) );
oa22f01  g5999 ( .o(n4308), .a(n5907), .b(n10294), .c(n5905), .d(n5570) );
na02f01  g6000 ( .o(n11488), .a(n7358), .b(_net_233) );
na02f01  g6001 ( .o(n11489), .a(n7352), .b(net_9664) );
ao22f01  g6002 ( .o(n11490), .a(n7357), .b(_net_10097), .c(n7353), .d(x5961) );
na04f01  g6003 ( .o(n4321), .a(n11490), .b(n11489), .c(n11488), .d(n7355_1) );
in01f01  g6004 ( .o(n11492), .a(net_10079) );
oa22f01  g6005 ( .o(n4326), .a(n6989_1), .b(n5618), .c(n6988), .d(n11492) );
no02f01  g6006 ( .o(n11494), .a(n9814), .b(_net_9296) );
na02f01  g6007 ( .o(n11495), .a(n9817), .b(n8809_1) );
oa22f01  g6008 ( .o(n4331), .a(n11495), .b(n11494), .c(n8817), .d(n7545) );
na02f01  g6009 ( .o(n11497), .a(n6038), .b(net_243) );
na02f01  g6010 ( .o(n11498), .a(n6037_1), .b(net_9872) );
ao22f01  g6011 ( .o(n11499), .a(n6044), .b(x5364), .c(n6042_1), .d(_net_10317) );
na04f01  g6012 ( .o(n4336), .a(n11499), .b(n11498), .c(n11497), .d(n6040) );
na03f01  g6013 ( .o(n11501), .a(n6068), .b(n5697), .c(_net_9512) );
ao12f01  g6014 ( .o(n11502), .a(_net_9421), .b(n6068), .c(_net_9512) );
no02f01  g6015 ( .o(n11503), .a(n11502), .b(n5697) );
ao22f01  g6016 ( .o(n11504), .a(n11503), .b(x2027), .c(n11502), .d(_net_9409) );
oa12f01  g6017 ( .o(n4341), .a(n11504), .b(n11501), .c(n10271) );
in01f01  g6018 ( .o(n11506), .a(_net_10255) );
no02f01  g6019 ( .o(n11507), .a(n6823), .b(n11506) );
in01f01  g6020 ( .o(n11508), .a(n6823) );
oa12f01  g6021 ( .o(n11509), .a(n6177_1), .b(n11508), .c(_net_10255) );
no02f01  g6022 ( .o(n11510), .a(n6842), .b(_net_10255) );
no03f01  g6023 ( .o(n11511), .a(n11510), .b(n6844), .c(n6846_1) );
ao12f01  g6024 ( .o(n11512), .a(n11511), .b(n6168), .c(_net_10255) );
oa12f01  g6025 ( .o(n4346), .a(n11512), .b(n11509), .c(n11507) );
na02f01  g6026 ( .o(n11514), .a(net_10194), .b(net_10180) );
ao22f01  g6027 ( .o(n11515), .a(net_10195), .b(net_10181), .c(net_10193), .d(net_10179) );
ao22f01  g6028 ( .o(n11516), .a(net_10189), .b(net_10176), .c(net_10192), .d(net_10179) );
ao22f01  g6029 ( .o(n11517), .a(net_10177), .b(net_10190), .c(net_10191), .d(net_10178) );
na04f01  g6030 ( .o(n4355), .a(n11517), .b(n11516), .c(n11515), .d(n11514) );
in01f01  g6031 ( .o(n11519), .a(n9679) );
in01f01  g6032 ( .o(n11520), .a(n9680) );
no02f01  g6033 ( .o(n11521), .a(n11520), .b(n9670) );
na03f01  g6034 ( .o(n11522), .a(n11521), .b(n11519), .c(n9673) );
in01f01  g6035 ( .o(n11523), .a(n11521) );
oa12f01  g6036 ( .o(n11524), .a(n11523), .b(n9679), .c(n9674) );
na02f01  g6037 ( .o(n4360), .a(n11524), .b(n11522) );
oa22f01  g6038 ( .o(n4372), .a(n5694), .b(n9579), .c(n5692), .d(n5609) );
na02f01  g6039 ( .o(n11527), .a(n6056), .b(net_236) );
na02f01  g6040 ( .o(n11528), .a(n6055), .b(net_9964) );
ao22f01  g6041 ( .o(n11529), .a(n6062_1), .b(x5790), .c(n6060), .d(_net_10415) );
na04f01  g6042 ( .o(n4377), .a(n11529), .b(n11528), .c(n11527), .d(n6058) );
ao12f01  g6043 ( .o(n11531), .a(n7530), .b(n6028_1), .c(n5994) );
oa12f01  g6044 ( .o(n4382), .a(n11531), .b(n6022), .c(n5990) );
in01f01  g6045 ( .o(n11533), .a(n5857) );
no03f01  g6046 ( .o(n11534), .a(n10356), .b(n11533), .c(n5884) );
in01f01  g6047 ( .o(n11535), .a(n8412) );
na02f01  g6048 ( .o(n11536), .a(net_9534), .b(n5489) );
no03f01  g6049 ( .o(n11537), .a(n11536), .b(n11535), .c(_net_9250) );
na02f01  g6050 ( .o(n11538), .a(_net_9503), .b(n8399_1) );
oa22f01  g6051 ( .o(n11539), .a(n11536), .b(n5871), .c(n11538), .d(n5891) );
no03f01  g6052 ( .o(n11540), .a(n11539), .b(n11537), .c(n11534) );
na03f01  g6053 ( .o(n11541), .a(n5880), .b(n5879), .c(net_9534) );
na02f01  g6054 ( .o(n11542), .a(n5891), .b(n5888_1) );
na03f01  g6055 ( .o(n11543), .a(n11542), .b(net_9534), .c(n8399_1) );
na03f01  g6056 ( .o(n4387), .a(n11543), .b(n11541), .c(n11540) );
oa22f01  g6057 ( .o(n4392), .a(n5694), .b(n5818), .c(n5692), .d(n5612) );
ao12f01  g6058 ( .o(n11546), .a(n5658), .b(n6532), .c(_net_259) );
ao22f01  g6059 ( .o(n11547), .a(n6535), .b(x4117), .c(n6534), .d(net_10019) );
na02f01  g6060 ( .o(n4397), .a(n11547), .b(n11546) );
na02f01  g6061 ( .o(n11549), .a(n8935), .b(_net_10327) );
na02f01  g6062 ( .o(n4405), .a(n11549), .b(n8937) );
oa22f01  g6063 ( .o(n11551), .a(n6600), .b(n6776), .c(n6563), .d(n8254) );
na02f01  g6064 ( .o(n11552), .a(n6584_1), .b(net_9770) );
na02f01  g6065 ( .o(n11553), .a(n6573), .b(net_9869) );
ao22f01  g6066 ( .o(n11554), .a(n6597), .b(_net_9735), .c(n6555), .d(net_9968) );
na03f01  g6067 ( .o(n11555), .a(n11554), .b(n11553), .c(n11552) );
no02f01  g6068 ( .o(n11556), .a(n11555), .b(n11551) );
in01f01  g6069 ( .o(n11557), .a(net_10000) );
oa22f01  g6070 ( .o(n11558), .a(n6966_1), .b(n5719_1), .c(n6959), .d(n11557) );
ao12f01  g6071 ( .o(n11559), .a(n11558), .b(n6585), .c(net_9703) );
ao22f01  g6072 ( .o(n11560), .a(n6582), .b(net_9901), .c(n6577), .d(net_9671) );
ao22f01  g6073 ( .o(n11561), .a(n6590), .b(_net_10032), .c(n6580), .d(net_9802) );
na04f01  g6074 ( .o(n4410), .a(n11561), .b(n11560), .c(n11559), .d(n11556) );
no02f01  g6075 ( .o(n11563), .a(n7375_1), .b(n7374) );
ao12f01  g6076 ( .o(n11564), .a(n7875), .b(n11563), .c(n7422) );
oa12f01  g6077 ( .o(n11565), .a(n11564), .b(n11563), .c(n7422) );
na02f01  g6078 ( .o(n11566), .a(n7444), .b(_net_10475) );
in01f01  g6079 ( .o(n11567), .a(n7444) );
ao12f01  g6080 ( .o(n11568), .a(n7451_1), .b(n11567), .c(n7373) );
ao22f01  g6081 ( .o(n11569), .a(n11568), .b(n11566), .c(n7453), .d(_net_10475) );
na02f01  g6082 ( .o(n4415), .a(n11569), .b(n11565) );
in01f01  g6083 ( .o(n11571), .a(n7596) );
in01f01  g6084 ( .o(n11572), .a(n7576) );
na02f01  g6085 ( .o(n11573), .a(n7584), .b(n11572) );
ao12f01  g6086 ( .o(n11574), .a(n11346), .b(n11573), .c(n11571) );
oa12f01  g6087 ( .o(n11575), .a(n11574), .b(n11573), .c(n11571) );
no02f01  g6088 ( .o(n11576), .a(n11345), .b(n7500) );
no02f01  g6089 ( .o(n11577), .a(n11345), .b(_net_9606) );
ao22f01  g6090 ( .o(n11578), .a(n11577), .b(_net_9602), .c(n11576), .d(net_102) );
na02f01  g6091 ( .o(n4420), .a(n11578), .b(n11575) );
no03f01  g6092 ( .o(n11580), .a(n7482), .b(n6485), .c(n6520) );
ao12f01  g6093 ( .o(n11581), .a(_net_9235), .b(n6490), .c(_net_9243) );
na02f01  g6094 ( .o(n11582), .a(n6476), .b(_net_9243) );
no03f01  g6095 ( .o(n11583), .a(n6497), .b(_net_9169), .c(n6520) );
ao12f01  g6096 ( .o(n11584), .a(n11583), .b(n6496), .c(_net_9243) );
na03f01  g6097 ( .o(n11585), .a(n11584), .b(n11582), .c(n11581) );
oa12f01  g6098 ( .o(n11586), .a(_net_9243), .b(n6492), .c(n6864) );
na02f01  g6099 ( .o(n11587), .a(n6471), .b(_net_9243) );
oa12f01  g6100 ( .o(n11588), .a(n11586), .b(n11587), .c(n7863) );
no03f01  g6101 ( .o(n11589), .a(n11588), .b(n11585), .c(n11580) );
no03f01  g6102 ( .o(n11590), .a(n6474_1), .b(n6520), .c(n6463) );
no03f01  g6103 ( .o(n11591), .a(n6861_1), .b(n6520), .c(n6511) );
ao12f01  g6104 ( .o(n11592), .a(n11587), .b(n7862_1), .c(n7852) );
no03f01  g6105 ( .o(n11593), .a(n11592), .b(n11591), .c(n11590) );
ao12f01  g6106 ( .o(n4425), .a(n6526_1), .b(n11593), .c(n11589) );
na02f01  g6107 ( .o(n11595), .a(n7937), .b(net_250) );
na02f01  g6108 ( .o(n11596), .a(n7936), .b(net_9780) );
ao22f01  g6109 ( .o(n11597), .a(n7943), .b(_net_10219), .c(n7942), .d(x4851) );
na04f01  g6110 ( .o(n4434), .a(n11597), .b(n11596), .c(n11595), .d(n7939) );
ao22f01  g6111 ( .o(n11599), .a(n5842), .b(net_9726), .c(n5841), .d(_net_167) );
na02f01  g6112 ( .o(n11600), .a(n5847), .b(net_10023) );
ao22f01  g6113 ( .o(n11601), .a(n5850), .b(net_9825), .c(n5849_1), .d(net_9924) );
na03f01  g6114 ( .o(n4439), .a(n11601), .b(n11600), .c(n11599) );
na02f01  g6115 ( .o(n11603), .a(n6038), .b(net_260) );
na02f01  g6116 ( .o(n11604), .a(n6037_1), .b(net_9889) );
ao22f01  g6117 ( .o(n11605), .a(n6044), .b(x4041), .c(n6042_1), .d(_net_10334) );
na04f01  g6118 ( .o(n4444), .a(n11605), .b(n11604), .c(n11603), .d(n6040) );
na02f01  g6119 ( .o(n11607), .a(n7358), .b(net_251) );
na02f01  g6120 ( .o(n11608), .a(n7352), .b(net_9682) );
ao22f01  g6121 ( .o(n11609), .a(n7357), .b(_net_10115), .c(n7353), .d(x4781) );
na04f01  g6122 ( .o(n4449), .a(n11609), .b(n11608), .c(n11607), .d(n7355_1) );
na02f01  g6123 ( .o(n11611), .a(n7353), .b(x5601) );
na02f01  g6124 ( .o(n11612), .a(n7352), .b(net_9670) );
ao22f01  g6125 ( .o(n11613), .a(n7358), .b(net_239), .c(n7357), .d(_net_10103) );
na04f01  g6126 ( .o(n4454), .a(n11613), .b(n11612), .c(n11611), .d(n7355_1) );
na02f01  g6127 ( .o(n11615), .a(n6760), .b(_net_10153) );
no02f01  g6128 ( .o(n11616), .a(n7782_1), .b(n7785) );
oa12f01  g6129 ( .o(n11617), .a(n6750), .b(n11616), .c(n8140_1) );
in01f01  g6130 ( .o(n11618), .a(n8127) );
na03f01  g6131 ( .o(n11619), .a(n8130_1), .b(n8128), .c(n11618) );
in01f01  g6132 ( .o(n11620), .a(n8128) );
oa12f01  g6133 ( .o(n11621), .a(n11620), .b(n8129), .c(n8127) );
na03f01  g6134 ( .o(n11622), .a(n11621), .b(n11619), .c(n10948) );
na03f01  g6135 ( .o(n4459), .a(n11622), .b(n11617), .c(n11615) );
ao22f01  g6136 ( .o(n11624), .a(n11503), .b(x1911), .c(n11502), .d(_net_9411) );
oa12f01  g6137 ( .o(n4468), .a(n11624), .b(n11501), .c(n8805) );
no02f01  g6138 ( .o(n11626), .a(n8269), .b(net_203) );
na02f01  g6139 ( .o(n11627), .a(n8272_1), .b(n573) );
oa22f01  g6140 ( .o(n4473), .a(n11627), .b(n11626), .c(n8280), .d(n8257) );
in01f01  g6141 ( .o(n11629), .a(net_10283) );
oa22f01  g6142 ( .o(n4482), .a(n9353), .b(n5609), .c(n9352), .d(n11629) );
in01f01  g6143 ( .o(n11631), .a(net_9540) );
no02f01  g6144 ( .o(n4487), .a(_net_9541), .b(n11631) );
in01f01  g6145 ( .o(n11633), .a(net_10300) );
na02f01  g6146 ( .o(n11634), .a(_net_9117), .b(net_10280) );
ao12f01  g6147 ( .o(n4496), .a(n5911), .b(n11634), .c(n11633) );
oa22f01  g6148 ( .o(n4501), .a(n9353), .b(n5597_1), .c(n9352), .d(n8610) );
ao12f01  g6149 ( .o(n11637), .a(n5658), .b(n6875_1), .c(net_258) );
ao22f01  g6150 ( .o(n11638), .a(n6878), .b(x4209), .c(n6877), .d(net_9919) );
na02f01  g6151 ( .o(n4506), .a(n11638), .b(n11637) );
ao22f01  g6152 ( .o(n11640), .a(n5842), .b(_net_9730), .c(n5841), .d(_net_171) );
na02f01  g6153 ( .o(n11641), .a(n5847), .b(_net_10027) );
ao22f01  g6154 ( .o(n11642), .a(n5850), .b(_net_9829), .c(n5849_1), .d(_net_9928) );
na03f01  g6155 ( .o(n4511), .a(n11642), .b(n11641), .c(n11640) );
in01f01  g6156 ( .o(n11644), .a(_net_10535) );
no03f01  g6157 ( .o(n4521), .a(n11644), .b(net_10537), .c(x1074) );
ao12f01  g6158 ( .o(n11646), .a(n5658), .b(n6875_1), .c(net_257) );
ao22f01  g6159 ( .o(n11647), .a(n6878), .b(x4285), .c(n6877), .d(net_9918) );
na02f01  g6160 ( .o(n4525), .a(n11647), .b(n11646) );
ao12f01  g6161 ( .o(n11649), .a(n5658), .b(n6532), .c(net_250) );
ao22f01  g6162 ( .o(n11650), .a(n6535), .b(x4851), .c(n6534), .d(net_10010) );
na02f01  g6163 ( .o(n4530), .a(n11650), .b(n11649) );
no02f01  g6164 ( .o(n4539), .a(n6164_1), .b(n8199) );
ao22f01  g6165 ( .o(n11653), .a(n5842), .b(net_9714), .c(n5841), .d(_net_154) );
na02f01  g6166 ( .o(n11654), .a(n5847), .b(net_10011) );
ao22f01  g6167 ( .o(n11655), .a(n5850), .b(net_9813), .c(n5849_1), .d(net_9912) );
na03f01  g6168 ( .o(n4544), .a(n11655), .b(n11654), .c(n11653) );
na04f01  g6169 ( .o(n11657), .a(n8778), .b(net_9605), .c(net_313), .d(net_9604) );
oa12f01  g6170 ( .o(n11658), .a(n11657), .b(n8776), .c(_net_9250) );
na02f01  g6171 ( .o(n11659), .a(n11658), .b(_net_9643) );
na03f01  g6172 ( .o(n11660), .a(n9494), .b(n7967_1), .c(_net_9637) );
oa12f01  g6173 ( .o(n4549), .a(n11659), .b(n11660), .c(n8745) );
ao12f01  g6174 ( .o(n11662), .a(n5658), .b(n7844), .c(net_247) );
ao22f01  g6175 ( .o(n11663), .a(n7847), .b(x5077), .c(n7846), .d(net_9809) );
na02f01  g6176 ( .o(n4554), .a(n11663), .b(n11662) );
na02f01  g6177 ( .o(n11665), .a(n7358), .b(_net_254) );
na02f01  g6178 ( .o(n11666), .a(n7352), .b(net_9685) );
ao22f01  g6179 ( .o(n11667), .a(n7357), .b(_net_10118), .c(n7353), .d(x4520) );
na04f01  g6180 ( .o(n4559), .a(n11667), .b(n11666), .c(n11665), .d(n7355_1) );
na02f01  g6181 ( .o(n11669), .a(n8936), .b(n7044_1) );
na02f01  g6182 ( .o(n11670), .a(n8937), .b(_net_10328) );
na02f01  g6183 ( .o(n4564), .a(n11670), .b(n11669) );
ao12f01  g6184 ( .o(n11672), .a(n5658), .b(n5678), .c(net_235) );
ao22f01  g6185 ( .o(n11673), .a(n5681_1), .b(x5850), .c(n5680), .d(net_9698) );
na02f01  g6186 ( .o(n4569), .a(n11673), .b(n11672) );
in01f01  g6187 ( .o(n11675), .a(net_9996) );
oa22f01  g6188 ( .o(n11676), .a(n6959), .b(n11675), .c(n6598), .d(n6720) );
in01f01  g6189 ( .o(n11677), .a(n6572) );
oa22f01  g6190 ( .o(n11678), .a(n6966_1), .b(n5710_1), .c(n11677), .d(n11243) );
no02f01  g6191 ( .o(n11679), .a(n11678), .b(n11676) );
oa22f01  g6192 ( .o(n11680), .a(n8046_1), .b(n8718), .c(n6563), .d(n8258) );
ao12f01  g6193 ( .o(n11681), .a(n11680), .b(n6564), .c(net_10077) );
ao22f01  g6194 ( .o(n11682), .a(n6584_1), .b(net_9766), .c(n6577), .d(net_9667) );
ao22f01  g6195 ( .o(n11683), .a(n6603), .b(net_10509), .c(n6585), .d(net_9699) );
oa12f01  g6196 ( .o(n11684), .a(n11683), .b(n8302), .c(n5909) );
ao22f01  g6197 ( .o(n11685), .a(n6590), .b(_net_10028), .c(n6580), .d(net_9798) );
ao22f01  g6198 ( .o(n11686), .a(n6599_1), .b(_net_9830), .c(n6555), .d(net_9964) );
ao22f01  g6199 ( .o(n11687), .a(n6592), .b(net_10194), .c(n6573), .d(net_9865) );
ao22f01  g6200 ( .o(n11688), .a(n8042), .b(net_10525), .c(n6582), .d(net_9897) );
na04f01  g6201 ( .o(n11689), .a(n11688), .b(n11687), .c(n11686), .d(n11685) );
no02f01  g6202 ( .o(n11690), .a(n11689), .b(n11684) );
na04f01  g6203 ( .o(n4574), .a(n11690), .b(n11682), .c(n11681), .d(n11679) );
na02f01  g6204 ( .o(n11692), .a(n8746), .b(_net_9572) );
ao12f01  g6205 ( .o(n4579), .a(n5658), .b(n11692), .c(n7958) );
na02f01  g6206 ( .o(n11694), .a(n9661), .b(n8142) );
no02f01  g6207 ( .o(n11695), .a(n11694), .b(n9660) );
no03f01  g6208 ( .o(n11696), .a(n11695), .b(n9657), .c(n6749) );
ao22f01  g6209 ( .o(n11697), .a(n6751), .b(_net_10114), .c(n6725), .d(_net_10115) );
no02f01  g6210 ( .o(n11698), .a(n11697), .b(_net_10141) );
ao22f01  g6211 ( .o(n11699), .a(n6714), .b(_net_10116), .c(_net_10117), .d(n6713_1) );
oa12f01  g6212 ( .o(n11700), .a(n11699), .b(n11697), .c(n7780) );
ao12f01  g6213 ( .o(n11701), .a(n6714), .b(_net_10117), .c(n6713_1) );
ao22f01  g6214 ( .o(n11702), .a(n11701), .b(n7772), .c(n7771), .d(_net_10143) );
oa12f01  g6215 ( .o(n11703), .a(n11702), .b(n11700), .c(n11698) );
oa22f01  g6216 ( .o(n11704), .a(_net_10147), .b(n7807), .c(n7808), .d(_net_10146) );
in01f01  g6217 ( .o(n11705), .a(n11704) );
ao22f01  g6218 ( .o(n11706), .a(_net_10118), .b(n6738_1), .c(_net_10119), .d(n10961) );
na03f01  g6219 ( .o(n11707), .a(n11706), .b(n11705), .c(n11703) );
oa22f01  g6220 ( .o(n11708), .a(n10982), .b(_net_10118), .c(n5747), .d(n6738_1) );
na02f01  g6221 ( .o(n11709), .a(n11708), .b(n11705) );
na03f01  g6222 ( .o(n11710), .a(n11705), .b(n7801_1), .c(_net_10145) );
ao12f01  g6223 ( .o(n11711), .a(n10965), .b(n10967), .c(_net_10121) );
ao22f01  g6224 ( .o(n11712), .a(n11711), .b(n7808), .c(_net_10147), .d(n7807) );
na04f01  g6225 ( .o(n11713), .a(n11712), .b(n11710), .c(n11709), .d(n11707) );
oa22f01  g6226 ( .o(n11714), .a(_net_10150), .b(n9363), .c(_net_10151), .d(n6667) );
oa22f01  g6227 ( .o(n11715), .a(n7761), .b(_net_10148), .c(_net_10149), .d(n7822) );
no02f01  g6228 ( .o(n11716), .a(n11715), .b(n11714) );
na02f01  g6229 ( .o(n11717), .a(n11716), .b(n11713) );
oa12f01  g6230 ( .o(n11718), .a(_net_10148), .b(_net_10149), .c(n7822) );
no03f01  g6231 ( .o(n11719), .a(n11718), .b(n11714), .c(_net_10122) );
no03f01  g6232 ( .o(n11720), .a(n11714), .b(n10949), .c(_net_10123) );
oa12f01  g6233 ( .o(n11721), .a(_net_10150), .b(_net_10151), .c(n6667) );
no02f01  g6234 ( .o(n11722), .a(n11721), .b(_net_10124) );
no03f01  g6235 ( .o(n11723), .a(_net_9752), .b(n6749), .c(n8248) );
oa12f01  g6236 ( .o(n11724), .a(n11723), .b(n11155), .c(_net_10125) );
no04f01  g6237 ( .o(n11725), .a(n11724), .b(n11722), .c(n11720), .d(n11719) );
ao12f01  g6238 ( .o(n11726), .a(n11696), .b(n11725), .c(n11717) );
no04f01  g6239 ( .o(n4589), .a(n11726), .b(net_10198), .c(_net_10197), .d(net_10199) );
ao22f01  g6240 ( .o(n11728), .a(n5842), .b(net_9682), .c(n5841), .d(_net_120) );
na02f01  g6241 ( .o(n11729), .a(n5847), .b(net_9979) );
ao22f01  g6242 ( .o(n11730), .a(n5850), .b(net_9781), .c(n5849_1), .d(net_9880) );
na03f01  g6243 ( .o(n4594), .a(n11730), .b(n11729), .c(n11728) );
oa22f01  g6244 ( .o(n4603), .a(n6989_1), .b(n5591), .c(n6988), .d(n10698) );
oa22f01  g6245 ( .o(n4608), .a(n7480_1), .b(n6163), .c(n7478), .d(n5582_1) );
in01f01  g6246 ( .o(n11734), .a(_net_9851) );
no02f01  g6247 ( .o(n11735), .a(n11734), .b(_net_9850) );
in01f01  g6248 ( .o(n11736), .a(n11735) );
no03f01  g6249 ( .o(n11737), .a(_net_10266), .b(_net_10268), .c(_net_10267) );
na03f01  g6250 ( .o(n11738), .a(n11737), .b(n6902), .c(n9185) );
no04f01  g6251 ( .o(n11739), .a(_net_10261), .b(_net_10263), .c(_net_10262), .d(_net_10264) );
na02f01  g6252 ( .o(n11740), .a(n11739), .b(n6903) );
no02f01  g6253 ( .o(n11741), .a(n11740), .b(n11738) );
no02f01  g6254 ( .o(n4613), .a(n11741), .b(n11736) );
na03f01  g6255 ( .o(n11743), .a(n7477), .b(x4520), .c(x6599) );
oa12f01  g6256 ( .o(n4618), .a(n11743), .b(n9831), .c(n10845) );
in01f01  g6257 ( .o(n11745), .a(_net_10202) );
ao12f01  g6258 ( .o(n11746), .a(n5658), .b(n6887), .c(x5961) );
oa12f01  g6259 ( .o(n4623), .a(n11746), .b(n6885_1), .c(n11745) );
no03f01  g6260 ( .o(n11748), .a(n9540), .b(n7966), .c(n8579) );
na03f01  g6261 ( .o(n11749), .a(n9542), .b(_net_9645), .c(_net_9641) );
na02f01  g6262 ( .o(n11750), .a(n9544), .b(_net_9645) );
ao12f01  g6263 ( .o(n11751), .a(n9546), .b(n8774), .c(n8579) );
no02f01  g6264 ( .o(n11752), .a(n8779), .b(n11145) );
no03f01  g6265 ( .o(n11753), .a(n9551), .b(n8781), .c(n9489) );
no04f01  g6266 ( .o(n11754), .a(n11753), .b(n11752), .c(n11751), .d(_net_9644) );
na03f01  g6267 ( .o(n11755), .a(n11754), .b(n11750), .c(n11749) );
oa12f01  g6268 ( .o(n11756), .a(x6599), .b(n11755), .c(n11748) );
no02f01  g6269 ( .o(n4632), .a(n11756), .b(n2827) );
no02f01  g6270 ( .o(n4637), .a(n10632), .b(n5688) );
na03f01  g6271 ( .o(n11759), .a(n7902_1), .b(net_9269), .c(net_9270) );
in01f01  g6272 ( .o(n11760), .a(net_9270) );
na03f01  g6273 ( .o(n11761), .a(n7899), .b(n10172), .c(n11760) );
na02f01  g6274 ( .o(n11762), .a(n11761), .b(n11759) );
na03f01  g6275 ( .o(n11763), .a(n7905), .b(net_9269), .c(n11760) );
na03f01  g6276 ( .o(n11764), .a(n7906_1), .b(n10172), .c(net_9270) );
na02f01  g6277 ( .o(n11765), .a(n11764), .b(n11763) );
no02f01  g6278 ( .o(n4642), .a(n11765), .b(n11762) );
ao12f01  g6279 ( .o(n11767), .a(n5658), .b(n6875_1), .c(net_246) );
ao22f01  g6280 ( .o(n11768), .a(n6878), .b(x5143), .c(n6877), .d(net_9907) );
na02f01  g6281 ( .o(n4654), .a(n11768), .b(n11767) );
oa22f01  g6282 ( .o(n4659), .a(n7756), .b(n6357), .c(n7755), .d(n6557) );
ao12f01  g6283 ( .o(n11771), .a(n5658), .b(n6052_1), .c(x4781) );
oa12f01  g6284 ( .o(n4664), .a(n11771), .b(n6048), .c(n8227_1) );
ao12f01  g6285 ( .o(n11773), .a(n5658), .b(n5678), .c(net_240) );
ao22f01  g6286 ( .o(n11774), .a(n5681_1), .b(x5548), .c(n5680), .d(net_9703) );
na02f01  g6287 ( .o(n4673), .a(n11774), .b(n11773) );
oa12f01  g6288 ( .o(n11776), .a(n9202), .b(n9195), .c(n10866) );
no02f01  g6289 ( .o(n11777), .a(n9206), .b(n9193) );
in01f01  g6290 ( .o(n11778), .a(n11777) );
na02f01  g6291 ( .o(n11779), .a(n11778), .b(n11776) );
in01f01  g6292 ( .o(n11780), .a(n11776) );
na02f01  g6293 ( .o(n11781), .a(n11777), .b(n11780) );
na02f01  g6294 ( .o(n4678), .a(n11781), .b(n11779) );
ao22f01  g6295 ( .o(n11783), .a(n11503), .b(x2214), .c(n11502), .d(_net_9406) );
oa12f01  g6296 ( .o(n4687), .a(n11783), .b(n11501), .c(n5737) );
in01f01  g6297 ( .o(n4696), .a(n9397) );
ao12f01  g6298 ( .o(n11786), .a(n5658), .b(n6532), .c(_net_255) );
ao22f01  g6299 ( .o(n11787), .a(n6535), .b(x4449), .c(n6534), .d(net_10015) );
na02f01  g6300 ( .o(n4705), .a(n11787), .b(n11786) );
ao22f01  g6301 ( .o(n11789), .a(n5842), .b(net_9737), .c(n5841), .d(_net_178) );
na02f01  g6302 ( .o(n11790), .a(n5847), .b(net_10034) );
ao22f01  g6303 ( .o(n11791), .a(n5850), .b(net_9836), .c(n5849_1), .d(net_9935) );
na03f01  g6304 ( .o(n4710), .a(n11791), .b(n11790), .c(n11789) );
in01f01  g6305 ( .o(n11793), .a(x3698) );
na02f01  g6306 ( .o(n11794), .a(_net_10488), .b(_net_10487) );
no02f01  g6307 ( .o(n11795), .a(n11794), .b(n9010) );
in01f01  g6308 ( .o(n11796), .a(_net_10489) );
no02f01  g6309 ( .o(n11797), .a(n9011), .b(n11796) );
no03f01  g6310 ( .o(n11798), .a(n11797), .b(n11795), .c(n11793) );
in01f01  g6311 ( .o(n11799), .a(_net_10512) );
ao12f01  g6312 ( .o(n11800), .a(n5658), .b(n11799), .c(_net_10511) );
na02f01  g6313 ( .o(n11801), .a(n11800), .b(x962) );
oa22f01  g6314 ( .o(n4715), .a(n11801), .b(n11798), .c(n11800), .d(n5658) );
in01f01  g6315 ( .o(n11803), .a(net_10185) );
oa22f01  g6316 ( .o(n4719), .a(n7956), .b(n5546), .c(n7955), .d(n11803) );
in01f01  g6317 ( .o(n11805), .a(net_10051) );
oa22f01  g6318 ( .o(n4729), .a(n9533), .b(n10282), .c(n9532), .d(n11805) );
no02f01  g6319 ( .o(n11807), .a(n10952), .b(n10951) );
ao12f01  g6320 ( .o(n11808), .a(n6746), .b(n11807), .c(n10975) );
oa12f01  g6321 ( .o(n11809), .a(n11808), .b(n11807), .c(n10975) );
na02f01  g6322 ( .o(n11810), .a(n10988), .b(n10950) );
no02f01  g6323 ( .o(n11811), .a(n10989), .b(n10398) );
ao22f01  g6324 ( .o(n11812), .a(n11811), .b(n11810), .c(n6760), .d(_net_10148) );
na02f01  g6325 ( .o(n4734), .a(n11812), .b(n11809) );
ao22f01  g6326 ( .o(n11814), .a(n5842), .b(net_9704), .c(n5841), .d(net_144) );
na02f01  g6327 ( .o(n11815), .a(n5847), .b(net_10001) );
ao22f01  g6328 ( .o(n11816), .a(n5850), .b(net_9803), .c(n5849_1), .d(net_9902) );
na03f01  g6329 ( .o(n4739), .a(n11816), .b(n11815), .c(n11814) );
in01f01  g6330 ( .o(n11818), .a(n7973) );
no04f01  g6331 ( .o(n4744), .a(n8748), .b(n7975), .c(n11818), .d(n8744) );
no02f01  g6332 ( .o(n11820), .a(n9404), .b(n8089) );
in01f01  g6333 ( .o(n11821), .a(n11820) );
na02f01  g6334 ( .o(n11822), .a(n11821), .b(n8085) );
no02f01  g6335 ( .o(n11823), .a(n11821), .b(n8085) );
in01f01  g6336 ( .o(n11824), .a(n11823) );
na02f01  g6337 ( .o(n11825), .a(n11824), .b(n11822) );
oa22f01  g6338 ( .o(n4749), .a(n11825), .b(n9397), .c(n9407), .d(n8085) );
oa12f01  g6339 ( .o(n4754), .a(n8110), .b(_net_9640), .c(_net_9639) );
in01f01  g6340 ( .o(n11828), .a(_net_231) );
oa12f01  g6341 ( .o(n11829), .a(x6599), .b(n5674), .c(n8687) );
na02f01  g6342 ( .o(n11830), .a(n8689), .b(net_10175) );
oa22f01  g6343 ( .o(n4759), .a(n11830), .b(n11828), .c(n11829), .d(n11475) );
ao12f01  g6344 ( .o(n11832), .a(n5658), .b(n5678), .c(_net_233) );
ao22f01  g6345 ( .o(n11833), .a(n5681_1), .b(x5961), .c(n5680), .d(net_9696) );
na02f01  g6346 ( .o(n4764), .a(n11833), .b(n11832) );
na02f01  g6347 ( .o(n11835), .a(n6776), .b(n6928) );
oa12f01  g6348 ( .o(n11836), .a(n11835), .b(n6929_1), .c(n6924_1) );
na02f01  g6349 ( .o(n11837), .a(n11836), .b(n6922) );
no02f01  g6350 ( .o(n11838), .a(n11837), .b(n6913) );
oa22f01  g6351 ( .o(n11839), .a(n11838), .b(n6930), .c(n11836), .d(n6928) );
no02f01  g6352 ( .o(n11840), .a(n9185), .b(n6773_1) );
no02f01  g6353 ( .o(n11841), .a(_net_10265), .b(_net_9835) );
no02f01  g6354 ( .o(n11842), .a(n11841), .b(n11840) );
ao12f01  g6355 ( .o(n11843), .a(n6933), .b(n11842), .c(n11839) );
oa12f01  g6356 ( .o(n11844), .a(n11843), .b(n11842), .c(n11839) );
na02f01  g6357 ( .o(n11845), .a(n6945), .b(_net_10265) );
ao12f01  g6358 ( .o(n11846), .a(n6846_1), .b(n6946), .c(n9185) );
ao22f01  g6359 ( .o(n11847), .a(n11846), .b(n11845), .c(n6168), .d(_net_10265) );
na02f01  g6360 ( .o(n4769), .a(n11847), .b(n11844) );
no02f01  g6361 ( .o(n11849), .a(n7660_1), .b(net_9617) );
no03f01  g6362 ( .o(n4774), .a(n11849), .b(n6545), .c(net_9613) );
ao12f01  g6363 ( .o(n11851), .a(n5658), .b(n6875_1), .c(net_235) );
ao22f01  g6364 ( .o(n11852), .a(n6878), .b(x5850), .c(n6877), .d(net_9896) );
na02f01  g6365 ( .o(n4779), .a(n11852), .b(n11851) );
na02f01  g6366 ( .o(n11854), .a(n6038), .b(net_253) );
na02f01  g6367 ( .o(n11855), .a(n6037_1), .b(net_9882) );
ao22f01  g6368 ( .o(n11856), .a(n6044), .b(x4587), .c(n6042_1), .d(_net_10327) );
na04f01  g6369 ( .o(n4788), .a(n11856), .b(n11855), .c(n11854), .d(n6040) );
na02f01  g6370 ( .o(n11858), .a(n11824), .b(n8086_1) );
no02f01  g6371 ( .o(n11859), .a(n11824), .b(n8086_1) );
in01f01  g6372 ( .o(n11860), .a(n11859) );
na02f01  g6373 ( .o(n11861), .a(n11860), .b(n11858) );
oa22f01  g6374 ( .o(n4797), .a(n11861), .b(n9397), .c(n9407), .d(n8086_1) );
na02f01  g6375 ( .o(n11863), .a(net_10285), .b(net_10299) );
ao22f01  g6376 ( .o(n11864), .a(net_10298), .b(net_10284), .c(net_10286), .d(net_10300) );
ao22f01  g6377 ( .o(n11865), .a(net_10281), .b(net_10294), .c(net_10297), .d(net_10284) );
ao22f01  g6378 ( .o(n11866), .a(net_10282), .b(net_10295), .c(net_10283), .d(net_10296) );
na04f01  g6379 ( .o(n4802), .a(n11866), .b(n11865), .c(n11864), .d(n11863) );
ao22f01  g6380 ( .o(n11868), .a(n5842), .b(net_9711), .c(n5841), .d(_net_151) );
na02f01  g6381 ( .o(n11869), .a(n5847), .b(net_10008) );
ao22f01  g6382 ( .o(n11870), .a(n5850), .b(net_9810), .c(n5849_1), .d(net_9909) );
na03f01  g6383 ( .o(n4807), .a(n11870), .b(n11869), .c(n11868) );
ao12f01  g6384 ( .o(n11872), .a(n5658), .b(n6160_1), .c(x4359) );
oa12f01  g6385 ( .o(n4812), .a(n11872), .b(n6159), .c(n7808) );
ao12f01  g6386 ( .o(n11874), .a(n5658), .b(n6875_1), .c(_net_259) );
ao22f01  g6387 ( .o(n11875), .a(n6878), .b(x4117), .c(n6877), .d(net_9920) );
na02f01  g6388 ( .o(n4817), .a(n11875), .b(n11874) );
na02f01  g6389 ( .o(n11877), .a(n7937), .b(net_257) );
na02f01  g6390 ( .o(n11878), .a(n7936), .b(net_9787) );
ao22f01  g6391 ( .o(n11879), .a(n7943), .b(_net_10226), .c(n7942), .d(x4285) );
na04f01  g6392 ( .o(n4822), .a(n11879), .b(n11878), .c(n11877), .d(n7939) );
oa12f01  g6393 ( .o(n11881), .a(x6599), .b(n6529), .c(n8687) );
na02f01  g6394 ( .o(n11882), .a(n8689), .b(net_10490) );
oa22f01  g6395 ( .o(n4827), .a(n11882), .b(n11828), .c(n11881), .d(n11479) );
in01f01  g6396 ( .o(n11884), .a(net_9936) );
oa22f01  g6397 ( .o(n4832), .a(n5694), .b(n11884), .c(n5692), .d(n5634) );
na02f01  g6398 ( .o(n11886), .a(n6056), .b(net_247) );
na02f01  g6399 ( .o(n11887), .a(n6055), .b(net_9975) );
ao22f01  g6400 ( .o(n11888), .a(n6062_1), .b(x5077), .c(n6060), .d(_net_10426) );
na04f01  g6401 ( .o(n4837), .a(n11888), .b(n11887), .c(n11886), .d(n6058) );
ao12f01  g6402 ( .o(n11890), .a(n5658), .b(n6532), .c(net_243) );
ao22f01  g6403 ( .o(n11891), .a(n6535), .b(x5364), .c(n6534), .d(net_10003) );
na02f01  g6404 ( .o(n4846), .a(n11891), .b(n11890) );
ao12f01  g6405 ( .o(n11893), .a(n5658), .b(n6160_1), .c(x4587) );
oa12f01  g6406 ( .o(n4851), .a(n11893), .b(n6159), .c(n7771) );
in01f01  g6407 ( .o(n11895), .a(net_9506) );
ao22f01  g6408 ( .o(n11896), .a(n5743), .b(x1660), .c(n5742), .d(_net_9415) );
oa12f01  g6409 ( .o(n4856), .a(n11896), .b(n5741), .c(n11895) );
na02f01  g6410 ( .o(n11898), .a(n7358), .b(net_252) );
na02f01  g6411 ( .o(n11899), .a(n7352), .b(net_9683) );
ao22f01  g6412 ( .o(n11900), .a(n7357), .b(_net_10116), .c(n7353), .d(x4694) );
na04f01  g6413 ( .o(n4866), .a(n11900), .b(n11899), .c(n11898), .d(n7355_1) );
na02f01  g6414 ( .o(n11902), .a(n1454), .b(n7991) );
in01f01  g6415 ( .o(n11903), .a(_net_9519) );
no02f01  g6416 ( .o(n11904), .a(n7995), .b(n11903) );
oa12f01  g6417 ( .o(n11905), .a(n7998), .b(n11904), .c(n9460) );
no02f01  g6418 ( .o(n11906), .a(n8002), .b(n11903) );
no02f01  g6419 ( .o(n11907), .a(n11906), .b(n5658) );
na03f01  g6420 ( .o(n4871), .a(n11907), .b(n11905), .c(n11902) );
in01f01  g6421 ( .o(n11909), .a(net_10286) );
oa22f01  g6422 ( .o(n4879), .a(n9353), .b(n5525), .c(n9352), .d(n11909) );
in01f01  g6423 ( .o(n11911), .a(net_10080) );
oa22f01  g6424 ( .o(n4884), .a(n6989_1), .b(n5606), .c(n6988), .d(n11911) );
na02f01  g6425 ( .o(n11913), .a(net_140), .b(net_149) );
na02f01  g6426 ( .o(n11914), .a(net_137), .b(net_145) );
no02f01  g6427 ( .o(n11915), .a(n11914), .b(n11913) );
na03f01  g6428 ( .o(n11916), .a(n11915), .b(net_135), .c(net_141) );
na04f01  g6429 ( .o(n11917), .a(net_134), .b(net_142), .c(net_146), .d(net_148) );
na04f01  g6430 ( .o(n11918), .a(net_139), .b(net_147), .c(net_150), .d(net_144) );
no02f01  g6431 ( .o(n11919), .a(n11918), .b(n11917) );
na04f01  g6432 ( .o(n11920), .a(n11919), .b(net_136), .c(net_138), .d(net_143) );
no02f01  g6433 ( .o(n4889), .a(n11920), .b(n11916) );
ao22f01  g6434 ( .o(n11922), .a(n9089), .b(_net_10339), .c(_net_10338), .d(n9087) );
no02f01  g6435 ( .o(n11923), .a(_net_10337), .b(n9128) );
ao22f01  g6436 ( .o(n11924), .a(n9129), .b(_net_8841), .c(_net_10337), .d(n9128) );
oa12f01  g6437 ( .o(n11925), .a(n11922), .b(n11924), .c(n11923) );
in01f01  g6438 ( .o(n11926), .a(_net_10339) );
in01f01  g6439 ( .o(n11927), .a(_net_10338) );
ao12f01  g6440 ( .o(n11928), .a(n9087), .b(n9089), .c(_net_10339) );
ao22f01  g6441 ( .o(n11929), .a(n11928), .b(n11927), .c(_net_10353), .d(n11926) );
ao22f01  g6442 ( .o(n11930), .a(n9110), .b(net_10342), .c(net_10343), .d(n9112) );
ao22f01  g6443 ( .o(n11931), .a(n9106), .b(_net_10340), .c(n9104), .d(_net_10341) );
na02f01  g6444 ( .o(n11932), .a(n11931), .b(n11930) );
ao12f01  g6445 ( .o(n11933), .a(n11932), .b(n11929), .c(n11925) );
in01f01  g6446 ( .o(n11934), .a(net_10345) );
oa12f01  g6447 ( .o(n11935), .a(_net_10358), .b(n11934), .c(_net_10359) );
oa22f01  g6448 ( .o(n11936), .a(n11935), .b(net_10344), .c(net_10345), .d(n9077) );
in01f01  g6449 ( .o(n11937), .a(_net_10360) );
ao22f01  g6450 ( .o(n11938), .a(n11937), .b(_net_10346), .c(n10140), .d(_net_10347) );
in01f01  g6451 ( .o(n11939), .a(_net_10347) );
oa12f01  g6452 ( .o(n11940), .a(_net_10360), .b(_net_10361), .c(n11939) );
oa22f01  g6453 ( .o(n11941), .a(n11940), .b(_net_10346), .c(n10140), .d(_net_10347) );
ao12f01  g6454 ( .o(n11942), .a(n11941), .b(n11938), .c(n11936) );
in01f01  g6455 ( .o(n11943), .a(_net_10341) );
oa12f01  g6456 ( .o(n11944), .a(_net_10354), .b(_net_10355), .c(n11943) );
oa22f01  g6457 ( .o(n11945), .a(n11944), .b(_net_10340), .c(n9104), .d(_net_10341) );
in01f01  g6458 ( .o(n11946), .a(net_10343) );
oa12f01  g6459 ( .o(n11947), .a(_net_10356), .b(n11946), .c(_net_10357) );
oa22f01  g6460 ( .o(n11948), .a(n11947), .b(net_10342), .c(net_10343), .d(n9112) );
ao12f01  g6461 ( .o(n11949), .a(n11948), .b(n11945), .c(n11930) );
na02f01  g6462 ( .o(n11950), .a(n11949), .b(n11942) );
in01f01  g6463 ( .o(n11951), .a(n11938) );
in01f01  g6464 ( .o(n11952), .a(net_10344) );
oa22f01  g6465 ( .o(n11953), .a(n11952), .b(_net_10358), .c(n11934), .d(_net_10359) );
oa12f01  g6466 ( .o(n11954), .a(n11942), .b(n11953), .c(n11951) );
oa12f01  g6467 ( .o(n4894), .a(n11954), .b(n11950), .c(n11933) );
ao22f01  g6468 ( .o(n11956), .a(n5842), .b(_net_9733), .c(n5841), .d(_net_174) );
na02f01  g6469 ( .o(n11957), .a(n5847), .b(_net_10030) );
ao22f01  g6470 ( .o(n11958), .a(n5850), .b(_net_9832), .c(n5849_1), .d(_net_9931) );
na03f01  g6471 ( .o(n4899), .a(n11958), .b(n11957), .c(n11956) );
oa22f01  g6472 ( .o(n4908), .a(n7756), .b(n5783), .c(n7755), .d(n10833) );
in01f01  g6473 ( .o(n11961), .a(_net_10112) );
ao12f01  g6474 ( .o(n11962), .a(n5658), .b(n6160_1), .c(x5003) );
oa12f01  g6475 ( .o(n4913), .a(n11962), .b(n6159), .c(n11961) );
in01f01  g6476 ( .o(n11964), .a(net_9836) );
oa22f01  g6477 ( .o(n4918), .a(n7480_1), .b(n11964), .c(n7478), .d(n5600) );
no03f01  g6478 ( .o(n11966), .a(n10776), .b(n10775), .c(_net_9204) );
no02f01  g6479 ( .o(n4923), .a(n11966), .b(n6686) );
no02f01  g6480 ( .o(n11968), .a(n9379), .b(n8334) );
no02f01  g6481 ( .o(n11969), .a(n9373), .b(_net_9326) );
no03f01  g6482 ( .o(n11970), .a(n11969), .b(n11968), .c(n10346) );
no02f01  g6483 ( .o(n11971), .a(n11969), .b(n11968) );
no02f01  g6484 ( .o(n11972), .a(n11971), .b(n10340) );
no02f01  g6485 ( .o(n11973), .a(_net_9323), .b(_net_9322) );
no02f01  g6486 ( .o(n11974), .a(n8759), .b(n8658) );
no02f01  g6487 ( .o(n11975), .a(n11974), .b(n11973) );
in01f01  g6488 ( .o(n11976), .a(n11975) );
no02f01  g6489 ( .o(n11977), .a(n11976), .b(n8639) );
no02f01  g6490 ( .o(n11978), .a(n11975), .b(_net_9319) );
no02f01  g6491 ( .o(n11979), .a(n11978), .b(n11977) );
in01f01  g6492 ( .o(n11980), .a(n11979) );
no03f01  g6493 ( .o(n11981), .a(n11980), .b(n11972), .c(n11970) );
no02f01  g6494 ( .o(n11982), .a(n11972), .b(n11970) );
no02f01  g6495 ( .o(n11983), .a(n11979), .b(n11982) );
no02f01  g6496 ( .o(n11984), .a(n11983), .b(n11981) );
no02f01  g6497 ( .o(n11985), .a(n11387), .b(net_9159) );
no02f01  g6498 ( .o(n11986), .a(n11386), .b(n8645) );
no02f01  g6499 ( .o(n11987), .a(n11986), .b(n11985) );
na02f01  g6500 ( .o(n11988), .a(n11987), .b(n11984) );
in01f01  g6501 ( .o(n11989), .a(n11984) );
in01f01  g6502 ( .o(n11990), .a(n11987) );
na02f01  g6503 ( .o(n11991), .a(n11990), .b(n11989) );
na03f01  g6504 ( .o(n11992), .a(n11991), .b(n11988), .c(n8638) );
ao12f01  g6505 ( .o(n11993), .a(n7883), .b(n8637), .c(_net_9311) );
na02f01  g6506 ( .o(n4932), .a(n11993), .b(n11992) );
no03f01  g6507 ( .o(n11995), .a(n10062), .b(n6491), .c(n6514) );
no02f01  g6508 ( .o(n4937), .a(n11995), .b(_net_9248) );
ao12f01  g6509 ( .o(n11997), .a(n5658), .b(n6532), .c(net_262) );
ao22f01  g6510 ( .o(n11998), .a(n6535), .b(x3889), .c(n6534), .d(net_10022) );
na02f01  g6511 ( .o(n4941), .a(n11998), .b(n11997) );
na02f01  g6512 ( .o(n12000), .a(n7353), .b(x5722) );
na02f01  g6513 ( .o(n12001), .a(n7352), .b(net_9668) );
ao22f01  g6514 ( .o(n12002), .a(n7358), .b(net_237), .c(n7357), .d(_net_10101) );
na04f01  g6515 ( .o(n4951), .a(n12002), .b(n12001), .c(n12000), .d(n7355_1) );
na02f01  g6516 ( .o(n12004), .a(n6056), .b(net_240) );
na02f01  g6517 ( .o(n12005), .a(n6055), .b(net_9968) );
ao22f01  g6518 ( .o(n12006), .a(n6062_1), .b(x5548), .c(n6060), .d(_net_10419) );
na04f01  g6519 ( .o(n4956), .a(n12006), .b(n12005), .c(n12004), .d(n6058) );
no02f01  g6520 ( .o(n12008), .a(n9105), .b(n9084) );
no03f01  g6521 ( .o(n12009), .a(n12008), .b(n9107), .c(n9101) );
oa12f01  g6522 ( .o(n12010), .a(n12008), .b(n9107), .c(n9101) );
na02f01  g6523 ( .o(n12011), .a(n12010), .b(n8183) );
no02f01  g6524 ( .o(n12012), .a(n9135), .b(n9106) );
oa12f01  g6525 ( .o(n12013), .a(n8200_1), .b(n12012), .c(_net_10355) );
ao12f01  g6526 ( .o(n12014), .a(n12013), .b(n12012), .c(_net_10355) );
ao12f01  g6527 ( .o(n12015), .a(n12014), .b(n8202), .c(_net_10355) );
oa12f01  g6528 ( .o(n4961), .a(n12015), .b(n12011), .c(n12009) );
no02f01  g6529 ( .o(n12017), .a(n10962), .b(n10958) );
no03f01  g6530 ( .o(n12018), .a(n12017), .b(n10955), .c(n6739) );
oa12f01  g6531 ( .o(n12019), .a(n12017), .b(n10955), .c(n6739) );
na02f01  g6532 ( .o(n12020), .a(n12019), .b(n10948) );
oa12f01  g6533 ( .o(n12021), .a(n6750), .b(n6758_1), .c(_net_10145) );
ao12f01  g6534 ( .o(n12022), .a(n12021), .b(n6758_1), .c(_net_10145) );
ao12f01  g6535 ( .o(n12023), .a(n12022), .b(n6760), .c(_net_10145) );
oa12f01  g6536 ( .o(n4971), .a(n12023), .b(n12020), .c(n12018) );
na02f01  g6537 ( .o(n12025), .a(n6038), .b(_net_255) );
na02f01  g6538 ( .o(n12026), .a(n6037_1), .b(net_9884) );
ao22f01  g6539 ( .o(n12027), .a(n6044), .b(x4449), .c(n6042_1), .d(_net_10329) );
na04f01  g6540 ( .o(n4980), .a(n12027), .b(n12026), .c(n12025), .d(n6040) );
in01f01  g6541 ( .o(n12029), .a(_net_10204) );
ao12f01  g6542 ( .o(n12030), .a(n5658), .b(n6887), .c(x5850) );
oa12f01  g6543 ( .o(n4985), .a(n12030), .b(n6885_1), .c(n12029) );
in01f01  g6544 ( .o(n12032), .a(_net_10418) );
ao12f01  g6545 ( .o(n12033), .a(n5658), .b(n6052_1), .c(x5601) );
oa12f01  g6546 ( .o(n4990), .a(n12033), .b(n6048), .c(n12032) );
oa12f01  g6547 ( .o(n12035), .a(n8917), .b(n8914), .c(n8918) );
oa12f01  g6548 ( .o(n12036), .a(n12035), .b(n8913), .c(n6014) );
in01f01  g6549 ( .o(n12037), .a(n8920) );
oa12f01  g6550 ( .o(n12038), .a(n12037), .b(n8909), .c(n8895) );
na03f01  g6551 ( .o(n12039), .a(n12038), .b(n12036), .c(net_9265) );
in01f01  g6552 ( .o(n12040), .a(net_9265) );
na02f01  g6553 ( .o(n12041), .a(n12038), .b(n12036) );
na02f01  g6554 ( .o(n12042), .a(n12041), .b(n12040) );
na02f01  g6555 ( .o(n4995), .a(n12042), .b(n12039) );
no03f01  g6556 ( .o(n12044), .a(n9540), .b(n7966), .c(n8783) );
na03f01  g6557 ( .o(n12045), .a(n9542), .b(_net_9646), .c(_net_9641) );
na02f01  g6558 ( .o(n12046), .a(n9495), .b(_net_9646) );
no02f01  g6559 ( .o(n12047), .a(n9546), .b(n8783) );
oa12f01  g6560 ( .o(n12048), .a(n8579), .b(n9791), .c(n8783) );
ao12f01  g6561 ( .o(n12049), .a(n12048), .b(n12047), .c(n8774) );
na03f01  g6562 ( .o(n12050), .a(n12049), .b(n12046), .c(n12045) );
oa12f01  g6563 ( .o(n12051), .a(x6599), .b(n12050), .c(n12044) );
no02f01  g6564 ( .o(n5000), .a(n12051), .b(n2827) );
na02f01  g6565 ( .o(n12053), .a(n7966), .b(_net_9637) );
oa22f01  g6566 ( .o(n5005), .a(n12053), .b(n7972_1), .c(n11657), .d(n11145) );
in01f01  g6567 ( .o(n12055), .a(net_10397) );
oa22f01  g6568 ( .o(n5010), .a(n10211), .b(n5552_1), .c(n10210), .d(n12055) );
ao22f01  g6569 ( .o(n12057), .a(n6714), .b(_net_10128), .c(n6713_1), .d(_net_10129) );
no02f01  g6570 ( .o(n12058), .a(n6725), .b(_net_10127) );
ao22f01  g6571 ( .o(n12059), .a(n6751), .b(_net_8845), .c(n6725), .d(_net_10127) );
oa12f01  g6572 ( .o(n12060), .a(n12057), .b(n12059), .c(n12058) );
in01f01  g6573 ( .o(n12061), .a(_net_10129) );
in01f01  g6574 ( .o(n12062), .a(_net_10128) );
ao12f01  g6575 ( .o(n12063), .a(n6714), .b(n6713_1), .c(_net_10129) );
ao22f01  g6576 ( .o(n12064), .a(n12063), .b(n12062), .c(_net_10143), .d(n12061) );
ao22f01  g6577 ( .o(n12065), .a(n10967), .b(net_10133), .c(n10965), .d(net_10132) );
ao22f01  g6578 ( .o(n12066), .a(_net_10131), .b(n10961), .c(_net_10130), .d(n6738_1) );
na02f01  g6579 ( .o(n12067), .a(n12066), .b(n12065) );
ao12f01  g6580 ( .o(n12068), .a(n12067), .b(n12064), .c(n12060) );
in01f01  g6581 ( .o(n12069), .a(net_10135) );
oa12f01  g6582 ( .o(n12070), .a(_net_10148), .b(_net_10149), .c(n12069) );
oa22f01  g6583 ( .o(n12071), .a(n12070), .b(net_10134), .c(n10949), .d(net_10135) );
in01f01  g6584 ( .o(n12072), .a(_net_10150) );
ao22f01  g6585 ( .o(n12073), .a(n12072), .b(_net_10136), .c(n11155), .d(_net_10137) );
in01f01  g6586 ( .o(n12074), .a(_net_10137) );
oa12f01  g6587 ( .o(n12075), .a(_net_10150), .b(_net_10151), .c(n12074) );
oa22f01  g6588 ( .o(n12076), .a(n12075), .b(_net_10136), .c(n11155), .d(_net_10137) );
ao12f01  g6589 ( .o(n12077), .a(n12076), .b(n12073), .c(n12071) );
in01f01  g6590 ( .o(n12078), .a(_net_10131) );
oa12f01  g6591 ( .o(n12079), .a(_net_10144), .b(n12078), .c(_net_10145) );
oa22f01  g6592 ( .o(n12080), .a(n12079), .b(_net_10130), .c(_net_10131), .d(n10961) );
in01f01  g6593 ( .o(n12081), .a(net_10133) );
oa12f01  g6594 ( .o(n12082), .a(_net_10146), .b(_net_10147), .c(n12081) );
oa22f01  g6595 ( .o(n12083), .a(n12082), .b(net_10132), .c(n10967), .d(net_10133) );
ao12f01  g6596 ( .o(n12084), .a(n12083), .b(n12080), .c(n12065) );
na02f01  g6597 ( .o(n12085), .a(n12084), .b(n12077) );
in01f01  g6598 ( .o(n12086), .a(n12073) );
in01f01  g6599 ( .o(n12087), .a(net_10134) );
oa22f01  g6600 ( .o(n12088), .a(n12087), .b(_net_10148), .c(_net_10149), .d(n12069) );
oa12f01  g6601 ( .o(n12089), .a(n12077), .b(n12088), .c(n12086) );
oa12f01  g6602 ( .o(n5015), .a(n12089), .b(n12085), .c(n12068) );
ao12f01  g6603 ( .o(n12091), .a(n5658), .b(n5774), .c(x4851) );
oa12f01  g6604 ( .o(n5020), .a(n12091), .b(n5770), .c(n3480) );
ao22f01  g6605 ( .o(n12093), .a(n8118), .b(x2890), .c(n8117), .d(_net_9395) );
oa12f01  g6606 ( .o(n5025), .a(n12093), .b(n8116_1), .c(n8805) );
ao12f01  g6607 ( .o(n12095), .a(n5658), .b(n7844), .c(_net_233) );
ao22f01  g6608 ( .o(n12096), .a(n7847), .b(x5961), .c(n7846), .d(net_9795) );
na02f01  g6609 ( .o(n5030), .a(n12096), .b(n12095) );
no03f01  g6610 ( .o(n12098), .a(_net_9242), .b(_net_9246), .c(_net_9245) );
na04f01  g6611 ( .o(n5035), .a(n12098), .b(n10421), .c(n10127), .d(n8454) );
no02f01  g6612 ( .o(n12100), .a(n7416), .b(n7406) );
in01f01  g6613 ( .o(n12101), .a(n12100) );
ao12f01  g6614 ( .o(n12102), .a(n7875), .b(n12101), .c(n7405) );
oa12f01  g6615 ( .o(n12103), .a(n12102), .b(n12101), .c(n7405) );
na02f01  g6616 ( .o(n12104), .a(n7437), .b(_net_10471) );
na02f01  g6617 ( .o(n12105), .a(n12104), .b(n7439) );
ao22f01  g6618 ( .o(n12106), .a(n12105), .b(n7450), .c(n7453), .d(_net_10471) );
na02f01  g6619 ( .o(n5043), .a(n12106), .b(n12103) );
in01f01  g6620 ( .o(n12108), .a(_net_10428) );
ao12f01  g6621 ( .o(n12109), .a(n5658), .b(n6052_1), .c(x4937) );
oa12f01  g6622 ( .o(n5048), .a(n12109), .b(n6048), .c(n12108) );
na03f01  g6623 ( .o(n12111), .a(n5746), .b(n7771), .c(n7772) );
na04f01  g6624 ( .o(n12112), .a(n7761), .b(n9363), .c(n6667), .d(n7822) );
no04f01  g6625 ( .o(n12113), .a(n12112), .b(n12111), .c(_net_10121), .d(_net_10120) );
no03f01  g6626 ( .o(n5057), .a(n12113), .b(_net_9752), .c(n8248) );
oa22f01  g6627 ( .o(n5062), .a(n8418), .b(n8718), .c(n8417), .d(n5537_1) );
in01f01  g6628 ( .o(n12116), .a(net_10089) );
oa22f01  g6629 ( .o(n5067), .a(n6989_1), .b(n5597_1), .c(n6988), .d(n12116) );
ao12f01  g6630 ( .o(n12118), .a(n5658), .b(n6532), .c(_net_233) );
ao22f01  g6631 ( .o(n12119), .a(n6535), .b(x5961), .c(n6534), .d(net_9993) );
na02f01  g6632 ( .o(n5072), .a(n12119), .b(n12118) );
na02f01  g6633 ( .o(n12121), .a(n7937), .b(net_235) );
na02f01  g6634 ( .o(n12122), .a(n7936), .b(net_9765) );
ao22f01  g6635 ( .o(n12123), .a(n7943), .b(_net_10204), .c(n7942), .d(x5850) );
na04f01  g6636 ( .o(n5077), .a(n12123), .b(n12122), .c(n12121), .d(n7939) );
in01f01  g6637 ( .o(n12125), .a(_net_9502) );
na02f01  g6638 ( .o(n5082), .a(n7989), .b(n12125) );
in01f01  g6639 ( .o(n12127), .a(net_9727) );
oa22f01  g6640 ( .o(n5091), .a(n7367), .b(n12127), .c(n7365_1), .d(n5513_1) );
na02f01  g6641 ( .o(n12129), .a(net_10495), .b(net_10509) );
ao22f01  g6642 ( .o(n12130), .a(net_10510), .b(net_10496), .c(net_10494), .d(net_10508) );
ao22f01  g6643 ( .o(n12131), .a(net_10504), .b(net_10491), .c(net_10507), .d(net_10494) );
ao22f01  g6644 ( .o(n12132), .a(net_10505), .b(net_10492), .c(net_10506), .d(net_10493) );
na04f01  g6645 ( .o(n5096), .a(n12132), .b(n12131), .c(n12130), .d(n12129) );
na02f01  g6646 ( .o(n12134), .a(n7937), .b(_net_232) );
na02f01  g6647 ( .o(n12135), .a(n7936), .b(net_9762) );
ao22f01  g6648 ( .o(n12136), .a(n7943), .b(_net_10201), .c(n7942), .d(x6028) );
na04f01  g6649 ( .o(n5105), .a(n12136), .b(n12135), .c(n12134), .d(n7939) );
na02f01  g6650 ( .o(n12138), .a(n7358), .b(_net_261) );
na02f01  g6651 ( .o(n12139), .a(n7352), .b(net_9692) );
ao22f01  g6652 ( .o(n12140), .a(n7357), .b(_net_10125), .c(n7353), .d(x3949) );
na04f01  g6653 ( .o(n5110), .a(n12140), .b(n12139), .c(n12138), .d(n7355_1) );
in01f01  g6654 ( .o(n12142), .a(n11400) );
no02f01  g6655 ( .o(n12143), .a(n8649), .b(_net_9318) );
no02f01  g6656 ( .o(n12144), .a(n8642), .b(n8758) );
no03f01  g6657 ( .o(n12145), .a(n12144), .b(n12143), .c(n11393) );
no02f01  g6658 ( .o(n12146), .a(n12144), .b(n12143) );
no02f01  g6659 ( .o(n12147), .a(n12146), .b(n11392) );
no03f01  g6660 ( .o(n12148), .a(n12147), .b(n12145), .c(n12142) );
no02f01  g6661 ( .o(n12149), .a(n12147), .b(n12145) );
no02f01  g6662 ( .o(n12150), .a(n12149), .b(n11400) );
no02f01  g6663 ( .o(n12151), .a(n12150), .b(n12148) );
na02f01  g6664 ( .o(n12152), .a(n12151), .b(n11987) );
in01f01  g6665 ( .o(n12153), .a(n12151) );
na02f01  g6666 ( .o(n12154), .a(n12153), .b(n11990) );
na03f01  g6667 ( .o(n12155), .a(n12154), .b(n12152), .c(n8638) );
ao12f01  g6668 ( .o(n12156), .a(n7883), .b(n8637), .c(_net_9326) );
na02f01  g6669 ( .o(n5115), .a(n12156), .b(n12155) );
in01f01  g6670 ( .o(n12158), .a(_net_10056) );
in01f01  g6671 ( .o(n12159), .a(_net_10057) );
na02f01  g6672 ( .o(n5120), .a(n12159), .b(n12158) );
oa22f01  g6673 ( .o(n5125), .a(n5694), .b(n5710_1), .c(n5692), .d(n5537_1) );
no02f01  g6674 ( .o(n12162), .a(n10314), .b(n10649) );
oa12f01  g6675 ( .o(n12163), .a(n7431), .b(n11330), .c(_net_10465) );
na02f01  g6676 ( .o(n12164), .a(n11337), .b(_net_10465) );
ao12f01  g6677 ( .o(n12165), .a(n7451_1), .b(n11338), .c(n10649) );
ao22f01  g6678 ( .o(n12166), .a(n12165), .b(n12164), .c(n7453), .d(_net_10465) );
oa12f01  g6679 ( .o(n5130), .a(n12166), .b(n12163), .c(n12162) );
na02f01  g6680 ( .o(n12168), .a(n6038), .b(_net_261) );
na02f01  g6681 ( .o(n12169), .a(n6037_1), .b(net_9890) );
ao22f01  g6682 ( .o(n12170), .a(n6044), .b(x3949), .c(n6042_1), .d(_net_10335) );
na04f01  g6683 ( .o(n5135), .a(n12170), .b(n12169), .c(n12168), .d(n6040) );
ao22f01  g6684 ( .o(n12172), .a(n8118), .b(x3133), .c(n8117), .d(_net_9391) );
oa12f01  g6685 ( .o(n5143), .a(n12172), .b(n8116_1), .c(n11895) );
ao12f01  g6686 ( .o(n12174), .a(n5658), .b(n5678), .c(net_238) );
ao22f01  g6687 ( .o(n12175), .a(n5681_1), .b(x5647), .c(n5680), .d(net_9701) );
na02f01  g6688 ( .o(n5152), .a(n12175), .b(n12174) );
oa22f01  g6689 ( .o(n5169), .a(n7367), .b(n6749), .c(n7365_1), .d(n5582_1) );
na02f01  g6690 ( .o(n12178), .a(n7353), .b(x5225) );
na02f01  g6691 ( .o(n12179), .a(n7352), .b(net_9676) );
ao22f01  g6692 ( .o(n12180), .a(n7358), .b(net_245), .c(n7357), .d(_net_10109) );
na04f01  g6693 ( .o(n5174), .a(n12180), .b(n12179), .c(n12178), .d(n7355_1) );
in01f01  g6694 ( .o(n12182), .a(n10389) );
no02f01  g6695 ( .o(n12183), .a(n12182), .b(n7820) );
no02f01  g6696 ( .o(n12184), .a(n10389), .b(_net_10161) );
oa12f01  g6697 ( .o(n12185), .a(n10948), .b(n12184), .c(n12183) );
no02f01  g6698 ( .o(n12186), .a(n10395), .b(n7820) );
ao12f01  g6699 ( .o(n12187), .a(_net_10161), .b(n10394), .c(n7763_1) );
no03f01  g6700 ( .o(n12188), .a(n12187), .b(n12186), .c(n10398) );
ao12f01  g6701 ( .o(n12189), .a(n12188), .b(n6760), .c(_net_10161) );
na02f01  g6702 ( .o(n5179), .a(n12189), .b(n12185) );
na02f01  g6703 ( .o(n12191), .a(n7453), .b(_net_10469) );
na02f01  g6704 ( .o(n12192), .a(n7434), .b(_net_10469) );
na02f01  g6705 ( .o(n12193), .a(n7435), .b(n7388) );
na03f01  g6706 ( .o(n12194), .a(n12193), .b(n12192), .c(n7450) );
oa12f01  g6707 ( .o(n12195), .a(n7403_1), .b(n7394_1), .c(n7390) );
in01f01  g6708 ( .o(n12196), .a(n7403_1) );
no02f01  g6709 ( .o(n12197), .a(n7394_1), .b(n7390) );
na02f01  g6710 ( .o(n12198), .a(n12197), .b(n12196) );
na03f01  g6711 ( .o(n12199), .a(n12198), .b(n12195), .c(n7431) );
na03f01  g6712 ( .o(n5184), .a(n12199), .b(n12194), .c(n12191) );
na02f01  g6713 ( .o(n12201), .a(_net_10325), .b(n3480) );
na02f01  g6714 ( .o(n12202), .a(n7027), .b(_net_10324) );
na02f01  g6715 ( .o(n5189), .a(n12202), .b(n12201) );
ao12f01  g6716 ( .o(n12204), .a(n5658), .b(n7844), .c(net_260) );
ao22f01  g6717 ( .o(n12205), .a(n7847), .b(x4041), .c(n7846), .d(net_9822) );
na02f01  g6718 ( .o(n5198), .a(n12205), .b(n12204) );
ao22f01  g6719 ( .o(n12207), .a(n5842), .b(net_9673), .c(n5841), .d(net_111) );
na02f01  g6720 ( .o(n12208), .a(n5847), .b(net_9970) );
ao22f01  g6721 ( .o(n12209), .a(n5850), .b(net_9772), .c(n5849_1), .d(net_9871) );
na03f01  g6722 ( .o(n5203), .a(n12209), .b(n12208), .c(n12207) );
na02f01  g6723 ( .o(n12211), .a(n9065), .b(n9200) );
na02f01  g6724 ( .o(n12212), .a(n9066), .b(_net_10223) );
na02f01  g6725 ( .o(n5208), .a(n12212), .b(n12211) );
ao22f01  g6726 ( .o(n12214), .a(n5743), .b(x1598), .c(n5742), .d(_net_9416) );
oa12f01  g6727 ( .o(n5217), .a(n12214), .b(n5741), .c(n5696) );
ao22f01  g6728 ( .o(n12216), .a(n6599_1), .b(_net_9827), .c(n6572), .d(net_10401) );
ao22f01  g6729 ( .o(n12217), .a(n8042), .b(net_10522), .c(n6580), .d(net_9795) );
ao22f01  g6730 ( .o(n12218), .a(n8047), .b(_net_10061), .c(n6562), .d(_net_199) );
oa12f01  g6731 ( .o(n12219), .a(n12218), .b(n8046_1), .c(n8733) );
na02f01  g6732 ( .o(n12220), .a(n6602), .b(net_9993) );
ao22f01  g6733 ( .o(n12221), .a(n8051_1), .b(net_10541), .c(n6564), .d(net_10074) );
na02f01  g6734 ( .o(n12222), .a(n12221), .b(n12220) );
no02f01  g6735 ( .o(n12223), .a(n12222), .b(n12219) );
ao22f01  g6736 ( .o(n12224), .a(n6605), .b(net_10296), .c(n6592), .d(net_10191) );
ao22f01  g6737 ( .o(n12225), .a(n6585), .b(net_9696), .c(n6573), .d(net_9862) );
na02f01  g6738 ( .o(n12226), .a(n12225), .b(n12224) );
ao22f01  g6739 ( .o(n12227), .a(n6606), .b(_net_9926), .c(n6555), .d(net_9961) );
ao22f01  g6740 ( .o(n12228), .a(n6603), .b(net_10506), .c(n6577), .d(net_9664) );
ao22f01  g6741 ( .o(n12229), .a(n6590), .b(_net_10025), .c(n6584_1), .d(net_9763) );
ao22f01  g6742 ( .o(n12230), .a(n6597), .b(_net_9728), .c(n6582), .d(net_9894) );
na04f01  g6743 ( .o(n12231), .a(n12230), .b(n12229), .c(n12228), .d(n12227) );
no02f01  g6744 ( .o(n12232), .a(n12231), .b(n12226) );
na04f01  g6745 ( .o(n5222), .a(n12232), .b(n12223), .c(n12217), .d(n12216) );
no02f01  g6746 ( .o(n12234), .a(n8277), .b(net_207) );
na02f01  g6747 ( .o(n12235), .a(n9450), .b(n573) );
oa22f01  g6748 ( .o(n5227), .a(n12235), .b(n12234), .c(n8280), .d(n9448) );
na02f01  g6749 ( .o(n12237), .a(n10713), .b(n6355) );
na02f01  g6750 ( .o(n12238), .a(net_210), .b(_net_9302) );
no02f01  g6751 ( .o(n12239), .a(net_211), .b(net_9303) );
no02f01  g6752 ( .o(n12240), .a(n9237), .b(n6362) );
no02f01  g6753 ( .o(n12241), .a(_net_9301), .b(net_209) );
no02f01  g6754 ( .o(n12242), .a(n6357), .b(n6557) );
oa22f01  g6755 ( .o(n12243), .a(n12242), .b(n12241), .c(n12240), .d(n12239) );
ao12f01  g6756 ( .o(n12244), .a(n12243), .b(n12238), .c(n12237) );
no02f01  g6757 ( .o(n12245), .a(net_9306), .b(net_214) );
no02f01  g6758 ( .o(n12246), .a(n6407), .b(n9518) );
no02f01  g6759 ( .o(n12247), .a(_net_193), .b(net_216) );
no02f01  g6760 ( .o(n12248), .a(n5783), .b(n10833) );
oa22f01  g6761 ( .o(n12249), .a(n12248), .b(n12247), .c(n12246), .d(n12245) );
no02f01  g6762 ( .o(n12250), .a(net_9307), .b(net_215) );
no02f01  g6763 ( .o(n12251), .a(n6373_1), .b(n9577) );
no02f01  g6764 ( .o(n12252), .a(net_212), .b(net_9304) );
in01f01  g6765 ( .o(n12253), .a(net_212) );
no02f01  g6766 ( .o(n12254), .a(n12253), .b(n6367) );
oa22f01  g6767 ( .o(n12255), .a(n12254), .b(n12252), .c(n12251), .d(n12250) );
no02f01  g6768 ( .o(n12256), .a(net_194), .b(net_217) );
no02f01  g6769 ( .o(n12257), .a(n5779), .b(n7753_1) );
no02f01  g6770 ( .o(n12258), .a(net_195), .b(net_218) );
no02f01  g6771 ( .o(n12259), .a(n5787_1), .b(n10818) );
oa22f01  g6772 ( .o(n12260), .a(n12259), .b(n12258), .c(n12257), .d(n12256) );
no02f01  g6773 ( .o(n12261), .a(net_219), .b(net_196) );
in01f01  g6774 ( .o(n12262), .a(net_219) );
no02f01  g6775 ( .o(n12263), .a(n12262), .b(n5791) );
no02f01  g6776 ( .o(n12264), .a(net_9305), .b(net_213) );
no02f01  g6777 ( .o(n12265), .a(n6387), .b(n8284) );
oa22f01  g6778 ( .o(n12266), .a(n12265), .b(n12264), .c(n12263), .d(n12261) );
no04f01  g6779 ( .o(n12267), .a(n12266), .b(n12260), .c(n12255), .d(n12249) );
na02f01  g6780 ( .o(n12268), .a(n12267), .b(n12244) );
no04f01  g6781 ( .o(n5232), .a(n12268), .b(n6461), .c(n5633), .d(n6354) );
ao12f01  g6782 ( .o(n12270), .a(n5658), .b(n6875_1), .c(net_253) );
ao22f01  g6783 ( .o(n12271), .a(n6878), .b(x4587), .c(n6877), .d(net_9914) );
na02f01  g6784 ( .o(n5237), .a(n12271), .b(n12270) );
no02f01  g6785 ( .o(n12273), .a(n9699), .b(n9698) );
no03f01  g6786 ( .o(n12274), .a(n12273), .b(n9717), .c(n9701) );
oa12f01  g6787 ( .o(n12275), .a(n12273), .b(n9717), .c(n9701) );
na02f01  g6788 ( .o(n12276), .a(n12275), .b(n7431) );
no02f01  g6789 ( .o(n12277), .a(n9731), .b(n9025) );
oa12f01  g6790 ( .o(n12278), .a(n7450), .b(n12277), .c(_net_10460) );
ao12f01  g6791 ( .o(n12279), .a(n12278), .b(n12277), .c(_net_10460) );
ao12f01  g6792 ( .o(n12280), .a(n12279), .b(n7453), .c(_net_10460) );
oa12f01  g6793 ( .o(n5242), .a(n12280), .b(n12276), .c(n12274) );
ao12f01  g6794 ( .o(n12282), .a(n5658), .b(n5678), .c(net_251) );
ao22f01  g6795 ( .o(n12283), .a(n5681_1), .b(x4781), .c(n5680), .d(net_9714) );
na02f01  g6796 ( .o(n5247), .a(n12283), .b(n12282) );
ao22f01  g6797 ( .o(n12285), .a(n5842), .b(net_9710), .c(n5841), .d(net_150) );
na02f01  g6798 ( .o(n12286), .a(n5847), .b(net_10007) );
ao22f01  g6799 ( .o(n12287), .a(n5850), .b(net_9809), .c(n5849_1), .d(net_9908) );
na03f01  g6800 ( .o(n5252), .a(n12287), .b(n12286), .c(n12285) );
na02f01  g6801 ( .o(n12289), .a(n7937), .b(net_238) );
na02f01  g6802 ( .o(n12290), .a(n7936), .b(net_9768) );
ao22f01  g6803 ( .o(n12291), .a(n7943), .b(_net_10207), .c(n7942), .d(x5647) );
na04f01  g6804 ( .o(n5257), .a(n12291), .b(n12290), .c(n12289), .d(n7939) );
ao22f01  g6805 ( .o(n12293), .a(n5842), .b(net_9722), .c(n5841), .d(_net_162) );
na02f01  g6806 ( .o(n12294), .a(n5847), .b(net_10019) );
ao22f01  g6807 ( .o(n12295), .a(n5850), .b(net_9821), .c(n5849_1), .d(net_9920) );
na03f01  g6808 ( .o(n5270), .a(n12295), .b(n12294), .c(n12293) );
no02f01  g6809 ( .o(n12297), .a(n7171), .b(n7093) );
no02f01  g6810 ( .o(n12298), .a(n7151), .b(n7091_1) );
no02f01  g6811 ( .o(n12299), .a(n12298), .b(n12297) );
no02f01  g6812 ( .o(n12300), .a(n12299), .b(n7315) );
na02f01  g6813 ( .o(n12301), .a(n12299), .b(n7315) );
na02f01  g6814 ( .o(n12302), .a(n12301), .b(n6148) );
ao12f01  g6815 ( .o(n12303), .a(n6131_1), .b(n6147), .c(net_9369) );
oa12f01  g6816 ( .o(n5275), .a(n12303), .b(n12302), .c(n12300) );
na02f01  g6817 ( .o(n12305), .a(n6020), .b(n5976) );
oa12f01  g6818 ( .o(n5283), .a(n12305), .b(n6020), .c(n5975) );
na02f01  g6819 ( .o(n12307), .a(n6349), .b(n6209) );
oa22f01  g6820 ( .o(n5288), .a(n12307), .b(n6348), .c(n6349), .d(n12040) );
na02f01  g6821 ( .o(n12309), .a(n6349), .b(n6336_1) );
oa22f01  g6822 ( .o(n5293), .a(n12309), .b(n6348), .c(n6349), .d(n8917) );
no03f01  g6823 ( .o(n5302), .a(n5929), .b(n8579), .c(n8578) );
ao22f01  g6824 ( .o(n12312), .a(n5842), .b(_net_9734), .c(n5841), .d(_net_175) );
na02f01  g6825 ( .o(n12313), .a(n5847), .b(_net_10031) );
ao22f01  g6826 ( .o(n12314), .a(n5850), .b(_net_9833), .c(n5849_1), .d(_net_9932) );
na03f01  g6827 ( .o(n5311), .a(n12314), .b(n12313), .c(n12312) );
ao12f01  g6828 ( .o(n12316), .a(n5658), .b(n6160_1), .c(x4041) );
oa12f01  g6829 ( .o(n5316), .a(n12316), .b(n6159), .c(n9363) );
in01f01  g6830 ( .o(n12318), .a(n7781) );
na03f01  g6831 ( .o(n12319), .a(n7787_1), .b(n7783), .c(n12318) );
oa12f01  g6832 ( .o(n12320), .a(n7784), .b(n7786), .c(n7781) );
na02f01  g6833 ( .o(n5321), .a(n12320), .b(n12319) );
na02f01  g6834 ( .o(n12322), .a(n6175), .b(n6829) );
no02f01  g6835 ( .o(n12323), .a(n6829), .b(_net_9827) );
oa12f01  g6836 ( .o(n12324), .a(n6177_1), .b(n12323), .c(n6789) );
na02f01  g6837 ( .o(n12325), .a(n6168), .b(_net_10245) );
na03f01  g6838 ( .o(n5326), .a(n12325), .b(n12324), .c(n12322) );
ao22f01  g6839 ( .o(n12327), .a(n5702), .b(x2648), .c(n5701), .d(_net_9399) );
oa12f01  g6840 ( .o(n5331), .a(n12327), .b(n5700_1), .c(n11895) );
na02f01  g6841 ( .o(n12329), .a(n6689_1), .b(n6671) );
na04f01  g6842 ( .o(n12330), .a(_net_9204), .b(_net_9207), .c(n6691), .d(net_9208) );
no04f01  g6843 ( .o(n5336), .a(n12330), .b(n12329), .c(n7647), .d(n6686) );
no02f01  g6844 ( .o(n12332), .a(n10300), .b(n10299) );
ao12f01  g6845 ( .o(n12333), .a(n7875), .b(n12332), .c(n10312) );
oa12f01  g6846 ( .o(n12334), .a(n12333), .b(n12332), .c(n10312) );
na02f01  g6847 ( .o(n12335), .a(n11334), .b(n10298) );
no02f01  g6848 ( .o(n12336), .a(n11335), .b(n7451_1) );
ao22f01  g6849 ( .o(n12337), .a(n12336), .b(n12335), .c(n7453), .d(_net_10463) );
na02f01  g6850 ( .o(n5341), .a(n12337), .b(n12334) );
in01f01  g6851 ( .o(n12339), .a(net_9837) );
oa22f01  g6852 ( .o(n5346), .a(n7480_1), .b(n12339), .c(n7478), .d(n5634) );
in01f01  g6853 ( .o(n12341), .a(net_10063) );
in01f01  g6854 ( .o(n12342), .a(_net_9661) );
ao12f01  g6855 ( .o(n5355), .a(n6155_1), .b(n12342), .c(n12341) );
na02f01  g6856 ( .o(n12344), .a(n7358), .b(net_235) );
na02f01  g6857 ( .o(n12345), .a(n7352), .b(net_9666) );
ao22f01  g6858 ( .o(n12346), .a(n7357), .b(_net_10099), .c(n7353), .d(x5850) );
na04f01  g6859 ( .o(n5360), .a(n12346), .b(n12345), .c(n12344), .d(n7355_1) );
no02f01  g6860 ( .o(n12348), .a(n8271), .b(net_204) );
na02f01  g6861 ( .o(n12349), .a(n8274), .b(n573) );
oa22f01  g6862 ( .o(n5365), .a(n12349), .b(n12348), .c(n8280), .d(n8256) );
ao12f01  g6863 ( .o(n12351), .a(n5658), .b(n7844), .c(_net_231) );
ao22f01  g6864 ( .o(n12352), .a(n7847), .b(x6102), .c(n7846), .d(net_9793) );
na02f01  g6865 ( .o(n5379), .a(n12352), .b(n12351) );
ao22f01  g6866 ( .o(n12354), .a(n5842), .b(net_9742), .c(n5841), .d(_net_182) );
na02f01  g6867 ( .o(n12355), .a(n5847), .b(net_10039) );
ao22f01  g6868 ( .o(n12356), .a(n5850), .b(net_9841), .c(n5849_1), .d(net_9940) );
na03f01  g6869 ( .o(n5384), .a(n12356), .b(n12355), .c(n12354) );
oa22f01  g6870 ( .o(n12358), .a(_net_10269), .b(n6178), .c(_net_8844), .d(n6183) );
na02f01  g6871 ( .o(n12359), .a(_net_10269), .b(n6178) );
oa22f01  g6872 ( .o(n12360), .a(n6904), .b(_net_10271), .c(_net_10270), .d(n6785) );
ao12f01  g6873 ( .o(n12361), .a(n12360), .b(n12359), .c(n12358) );
in01f01  g6874 ( .o(n12362), .a(_net_10271) );
oa12f01  g6875 ( .o(n12363), .a(_net_10270), .b(n6904), .c(_net_10271) );
oa22f01  g6876 ( .o(n12364), .a(n12363), .b(_net_9829), .c(_net_9830), .d(n12362) );
no02f01  g6877 ( .o(n12365), .a(n12364), .b(n12361) );
oa22f01  g6878 ( .o(n12366), .a(n6799), .b(net_10274), .c(net_10275), .d(n6776) );
oa22f01  g6879 ( .o(n12367), .a(_net_10272), .b(n6778_1), .c(n6801_1), .d(_net_10273) );
no03f01  g6880 ( .o(n12368), .a(n12367), .b(n12366), .c(n12365) );
in01f01  g6881 ( .o(n12369), .a(_net_10273) );
in01f01  g6882 ( .o(n12370), .a(_net_10272) );
ao12f01  g6883 ( .o(n12371), .a(n12370), .b(_net_9832), .c(n12369) );
ao22f01  g6884 ( .o(n12372), .a(n12371), .b(n6778_1), .c(n6801_1), .d(_net_10273) );
oa12f01  g6885 ( .o(n12373), .a(net_10274), .b(net_10275), .c(n6776) );
no02f01  g6886 ( .o(n12374), .a(n12373), .b(_net_9833) );
ao12f01  g6887 ( .o(n12375), .a(n12374), .b(net_10275), .c(n6776) );
oa12f01  g6888 ( .o(n12376), .a(n12375), .b(n12372), .c(n12366) );
oa22f01  g6889 ( .o(n12377), .a(n12376), .b(n12368), .c(_net_10276), .d(n6773_1) );
na02f01  g6890 ( .o(n12378), .a(_net_10276), .b(n6773_1) );
no03f01  g6891 ( .o(n12379), .a(net_8816), .b(net_8837), .c(_net_8817) );
na03f01  g6892 ( .o(n5389), .a(n12379), .b(n12378), .c(n12377) );
na02f01  g6893 ( .o(n12381), .a(n6760), .b(_net_10141) );
na02f01  g6894 ( .o(n12382), .a(n6751), .b(n6725) );
na03f01  g6895 ( .o(n12383), .a(n12382), .b(n6753_1), .c(n6750) );
in01f01  g6896 ( .o(n12384), .a(n6728_1) );
no02f01  g6897 ( .o(n12385), .a(n6730), .b(n6726) );
na02f01  g6898 ( .o(n12386), .a(n12385), .b(n12384) );
oa12f01  g6899 ( .o(n12387), .a(n6728_1), .b(n6730), .c(n6726) );
na03f01  g6900 ( .o(n12388), .a(n12387), .b(n12386), .c(n10948) );
na03f01  g6901 ( .o(n5394), .a(n12388), .b(n12383), .c(n12381) );
ao22f01  g6902 ( .o(n12390), .a(n5842), .b(net_9688), .c(n5841), .d(_net_126) );
na02f01  g6903 ( .o(n12391), .a(n5847), .b(net_9985) );
ao22f01  g6904 ( .o(n12392), .a(n5850), .b(net_9787), .c(n5849_1), .d(net_9886) );
na03f01  g6905 ( .o(n5399), .a(n12392), .b(n12391), .c(n12390) );
ao12f01  g6906 ( .o(n12394), .a(n5658), .b(n6160_1), .c(x4449) );
oa12f01  g6907 ( .o(n5412), .a(n12394), .b(n6159), .c(n7801_1) );
na02f01  g6908 ( .o(n12396), .a(n7243), .b(n7100_1) );
na02f01  g6909 ( .o(n12397), .a(n7236), .b(n7099) );
na03f01  g6910 ( .o(n12398), .a(n12397), .b(n12396), .c(n6148) );
ao12f01  g6911 ( .o(n12399), .a(n6131_1), .b(n6147), .c(net_9365) );
na02f01  g6912 ( .o(n5417), .a(n12399), .b(n12398) );
no02f01  g6913 ( .o(n12401), .a(_net_10476), .b(n9043) );
no02f01  g6914 ( .o(n12402), .a(n7371), .b(_net_10438) );
in01f01  g6915 ( .o(n12403), .a(n12402) );
no02f01  g6916 ( .o(n12404), .a(n9044), .b(_net_10475) );
ao12f01  g6917 ( .o(n12405), .a(n12401), .b(n12404), .c(n12403) );
in01f01  g6918 ( .o(n12406), .a(n12405) );
no02f01  g6919 ( .o(n12407), .a(_net_10437), .b(n7373) );
no02f01  g6920 ( .o(n12408), .a(n7377), .b(_net_10436) );
in01f01  g6921 ( .o(n12409), .a(n8239) );
na02f01  g6922 ( .o(n12410), .a(n12409), .b(n8237) );
no02f01  g6923 ( .o(n12411), .a(n8239), .b(n8215) );
no02f01  g6924 ( .o(n12412), .a(_net_10474), .b(n9027) );
no02f01  g6925 ( .o(n12413), .a(n12412), .b(n8241) );
ao12f01  g6926 ( .o(n12414), .a(n12413), .b(n12408), .c(n9027) );
no02f01  g6927 ( .o(n12415), .a(n12414), .b(n12411) );
ao12f01  g6928 ( .o(n12416), .a(n12408), .b(n12415), .c(n12410) );
na02f01  g6929 ( .o(n12417), .a(n12414), .b(n7377) );
in01f01  g6930 ( .o(n12418), .a(n12417) );
no02f01  g6931 ( .o(n12419), .a(n12418), .b(n12416) );
no02f01  g6932 ( .o(n12420), .a(n12419), .b(n12407) );
na02f01  g6933 ( .o(n12421), .a(n12420), .b(n12403) );
in01f01  g6934 ( .o(n12422), .a(n12421) );
no02f01  g6935 ( .o(n12423), .a(n7370_1), .b(_net_10439) );
no02f01  g6936 ( .o(n12424), .a(_net_10477), .b(n9041) );
no02f01  g6937 ( .o(n12425), .a(n12424), .b(n12423) );
in01f01  g6938 ( .o(n12426), .a(n12425) );
oa12f01  g6939 ( .o(n12427), .a(n12426), .b(n12422), .c(n12406) );
na03f01  g6940 ( .o(n12428), .a(n12425), .b(n12421), .c(n12405) );
na02f01  g6941 ( .o(n5422), .a(n12428), .b(n12427) );
in01f01  g6942 ( .o(n12430), .a(n8533) );
na02f01  g6943 ( .o(n12431), .a(n10385), .b(n12430) );
no02f01  g6944 ( .o(n12432), .a(n12431), .b(n10383) );
no02f01  g6945 ( .o(n12433), .a(n10380), .b(n10378) );
in01f01  g6946 ( .o(n12434), .a(n12433) );
ao12f01  g6947 ( .o(n12435), .a(n6746), .b(n12434), .c(n12432) );
oa12f01  g6948 ( .o(n12436), .a(n12435), .b(n12434), .c(n12432) );
in01f01  g6949 ( .o(n12437), .a(n10394) );
na02f01  g6950 ( .o(n12438), .a(n8541), .b(_net_10159) );
na02f01  g6951 ( .o(n12439), .a(n12438), .b(n12437) );
ao22f01  g6952 ( .o(n12440), .a(n12439), .b(n6750), .c(n6760), .d(_net_10159) );
na02f01  g6953 ( .o(n5427), .a(n12440), .b(n12436) );
no02f01  g6954 ( .o(n12442), .a(n9122), .b(n11937) );
oa12f01  g6955 ( .o(n12443), .a(n8183), .b(n9123), .c(_net_10360) );
na02f01  g6956 ( .o(n12444), .a(n9143), .b(n11937) );
no02f01  g6957 ( .o(n12445), .a(n10145), .b(n9144) );
ao22f01  g6958 ( .o(n12446), .a(n12445), .b(n12444), .c(n8202), .d(_net_10360) );
oa12f01  g6959 ( .o(n5436), .a(n12446), .b(n12443), .c(n12442) );
no02f01  g6960 ( .o(n12448), .a(n6026), .b(n7593) );
ao12f01  g6961 ( .o(n12449), .a(n12448), .b(n6028_1), .c(n8841) );
oa12f01  g6962 ( .o(n5441), .a(n12449), .b(n6022), .c(n7592) );
ao12f01  g6963 ( .o(n12451), .a(n5658), .b(n5678), .c(net_242) );
ao22f01  g6964 ( .o(n12452), .a(n5681_1), .b(x5427), .c(n5680), .d(net_9705) );
na02f01  g6965 ( .o(n5454), .a(n12452), .b(n12451) );
no02f01  g6966 ( .o(n12454), .a(n9323), .b(n9322) );
ao12f01  g6967 ( .o(n12455), .a(n8184), .b(n12454), .c(n9329) );
oa12f01  g6968 ( .o(n12456), .a(n12455), .b(n12454), .c(n9329) );
na02f01  g6969 ( .o(n12457), .a(n9267), .b(_net_10370) );
ao12f01  g6970 ( .o(n12458), .a(n9144), .b(n9268), .c(n7003_1) );
ao22f01  g6971 ( .o(n12459), .a(n12458), .b(n12457), .c(n8202), .d(_net_10370) );
na02f01  g6972 ( .o(n5459), .a(n12459), .b(n12456) );
ao22f01  g6973 ( .o(n12461), .a(n11503), .b(x2165), .c(n11502), .d(_net_9407) );
oa12f01  g6974 ( .o(n5464), .a(n12461), .b(n11501), .c(n11895) );
oa22f01  g6975 ( .o(n12463), .a(n6565), .b(n10698), .c(n6563), .d(n10713) );
ao12f01  g6976 ( .o(n12464), .a(n12463), .b(n6555), .c(net_9976) );
ao22f01  g6977 ( .o(n12465), .a(n6573), .b(net_9877), .c(n6572), .d(net_10393) );
ao22f01  g6978 ( .o(n12466), .a(n6580), .b(net_9810), .c(n6577), .d(net_9679) );
na02f01  g6979 ( .o(n12467), .a(n6584_1), .b(net_9778) );
ao22f01  g6980 ( .o(n12468), .a(n6599_1), .b(net_9841), .c(n6582), .d(net_9909) );
na02f01  g6981 ( .o(n12469), .a(n12468), .b(n12467) );
ao22f01  g6982 ( .o(n12470), .a(n6592), .b(net_10183), .c(n6590), .d(net_10039) );
ao22f01  g6983 ( .o(n12471), .a(n6597), .b(net_9742), .c(n6585), .d(net_9711) );
ao22f01  g6984 ( .o(n12472), .a(n6603), .b(net_10498), .c(n6602), .d(net_10008) );
ao22f01  g6985 ( .o(n12473), .a(n6606), .b(net_9940), .c(n6605), .d(net_10288) );
na04f01  g6986 ( .o(n12474), .a(n12473), .b(n12472), .c(n12471), .d(n12470) );
no02f01  g6987 ( .o(n12475), .a(n12474), .b(n12469) );
na04f01  g6988 ( .o(n5469), .a(n12475), .b(n12466), .c(n12465), .d(n12464) );
in01f01  g6989 ( .o(n12477), .a(net_10402) );
na02f01  g6990 ( .o(n12478), .a(n9799), .b(net_10385) );
ao12f01  g6991 ( .o(n5481), .a(n11245), .b(n12478), .c(n12477) );
na03f01  g6992 ( .o(n12480), .a(_net_10325), .b(_net_10324), .c(_net_10326) );
na02f01  g6993 ( .o(n5486), .a(n12480), .b(n8935) );
in01f01  g6994 ( .o(n12482), .a(net_9260) );
na02f01  g6995 ( .o(n12483), .a(n6349), .b(n6230) );
oa22f01  g6996 ( .o(n5491), .a(n12483), .b(n6348), .c(n6349), .d(n12482) );
oa22f01  g6997 ( .o(n5500), .a(n7367), .b(n6727), .c(n7365_1), .d(n5621) );
na02f01  g6998 ( .o(n12486), .a(n6056), .b(_net_261) );
na02f01  g6999 ( .o(n12487), .a(n6055), .b(net_9989) );
ao22f01  g7000 ( .o(n12488), .a(n6062_1), .b(x3949), .c(n6060), .d(_net_10440) );
na04f01  g7001 ( .o(n5513), .a(n12488), .b(n12487), .c(n12486), .d(n6058) );
no04f01  g7002 ( .o(n12490), .a(net_9576), .b(net_9577), .c(_net_9581), .d(net_9583) );
na02f01  g7003 ( .o(n12491), .a(n12490), .b(n9883) );
na04f01  g7004 ( .o(n12492), .a(n9882), .b(n9847), .c(n9843), .d(n9876) );
na04f01  g7005 ( .o(n12493), .a(n9869), .b(n9846), .c(n9863), .d(n9861) );
no03f01  g7006 ( .o(n5518), .a(n12493), .b(n12492), .c(n12491) );
in01f01  g7007 ( .o(n12495), .a(_net_10305) );
ao12f01  g7008 ( .o(n12496), .a(n5658), .b(n5774), .c(x6102) );
oa12f01  g7009 ( .o(n5523), .a(n12496), .b(n5770), .c(n12495) );
na03f01  g7010 ( .o(n12498), .a(n8776), .b(n8399_1), .c(_net_9643) );
oa12f01  g7011 ( .o(n5528), .a(n12498), .b(n8751), .c(n7973) );
no02f01  g7012 ( .o(n12500), .a(n6561_1), .b(n11210) );
ao22f01  g7013 ( .o(n12501), .a(n12500), .b(n6558), .c(n6585), .d(net_9725) );
ao22f01  g7014 ( .o(n12502), .a(n6599_1), .b(net_9855), .c(n6584_1), .d(net_9792) );
ao22f01  g7015 ( .o(n12503), .a(n6573), .b(net_9891), .c(n6555), .d(net_9990) );
na02f01  g7016 ( .o(n12504), .a(n6582), .b(net_9923) );
ao22f01  g7017 ( .o(n12505), .a(n6580), .b(net_9824), .c(n6577), .d(net_9693) );
na02f01  g7018 ( .o(n12506), .a(n12505), .b(n12504) );
in01f01  g7019 ( .o(n12507), .a(net_9756) );
oa22f01  g7020 ( .o(n12508), .a(n6966_1), .b(n8685), .c(n6598), .d(n12507) );
in01f01  g7021 ( .o(n12509), .a(net_10022) );
in01f01  g7022 ( .o(n12510), .a(net_10053) );
oa22f01  g7023 ( .o(n12511), .a(n6959), .b(n12509), .c(n6591), .d(n12510) );
no03f01  g7024 ( .o(n12512), .a(n12511), .b(n12508), .c(n12506) );
na04f01  g7025 ( .o(n5533), .a(n12512), .b(n12503), .c(n12502), .d(n12501) );
ao12f01  g7026 ( .o(n12514), .a(n6921), .b(n9437), .c(n6915) );
in01f01  g7027 ( .o(n12515), .a(n12514) );
no02f01  g7028 ( .o(n12516), .a(n6924_1), .b(n6911) );
ao12f01  g7029 ( .o(n12517), .a(n6933), .b(n12516), .c(n12515) );
oa12f01  g7030 ( .o(n12518), .a(n12517), .b(n12516), .c(n12515) );
na02f01  g7031 ( .o(n12519), .a(n6942), .b(_net_10263) );
na02f01  g7032 ( .o(n12520), .a(n12519), .b(n6944_1) );
ao22f01  g7033 ( .o(n12521), .a(n12520), .b(n6175), .c(n6168), .d(_net_10263) );
na02f01  g7034 ( .o(n5537), .a(n12521), .b(n12518) );
ao12f01  g7035 ( .o(n12523), .a(n5658), .b(n6052_1), .c(x4117) );
oa12f01  g7036 ( .o(n5542), .a(n12523), .b(n6048), .c(n9043) );
ao22f01  g7037 ( .o(n12525), .a(n8118), .b(x3022), .c(n8117), .d(_net_9393) );
oa12f01  g7038 ( .o(n5547), .a(n12525), .b(n8116_1), .c(n10271) );
ao22f01  g7039 ( .o(n12527), .a(n5842), .b(_net_9740), .c(n5841), .d(_net_180) );
na02f01  g7040 ( .o(n12528), .a(n5847), .b(_net_10037) );
ao22f01  g7041 ( .o(n12529), .a(n5850), .b(_net_9839), .c(n5849_1), .d(_net_9938) );
na03f01  g7042 ( .o(n5552), .a(n12529), .b(n12528), .c(n12527) );
in01f01  g7043 ( .o(n12531), .a(net_9854) );
oa12f01  g7044 ( .o(n12532), .a(x6599), .b(n7841), .c(n8687) );
na02f01  g7045 ( .o(n12533), .a(n8689), .b(net_10280) );
oa22f01  g7046 ( .o(n5557), .a(n12533), .b(n11828), .c(n12532), .d(n12531) );
na02f01  g7047 ( .o(n12535), .a(n8695), .b(net_9159) );
oa12f01  g7048 ( .o(n5562), .a(n12535), .b(n8695), .c(n5783) );
in01f01  g7049 ( .o(n12537), .a(n9100) );
no02f01  g7050 ( .o(n12538), .a(n9107), .b(n9086) );
ao12f01  g7051 ( .o(n12539), .a(n8184), .b(n12538), .c(n12537) );
oa12f01  g7052 ( .o(n12540), .a(n12539), .b(n12538), .c(n12537) );
no02f01  g7053 ( .o(n12541), .a(n9134), .b(_net_10354) );
no02f01  g7054 ( .o(n12542), .a(n12541), .b(n12012) );
ao22f01  g7055 ( .o(n12543), .a(n12542), .b(n8200_1), .c(n8202), .d(_net_10354) );
na02f01  g7056 ( .o(n5567), .a(n12543), .b(n12540) );
no02f01  g7057 ( .o(n12545), .a(net_9615), .b(net_9614) );
no03f01  g7058 ( .o(n5572), .a(n12545), .b(n6543), .c(net_9613) );
na02f01  g7059 ( .o(n12547), .a(n6020), .b(n6617) );
oa12f01  g7060 ( .o(n5577), .a(n12547), .b(n6020), .c(n8468) );
in01f01  g7061 ( .o(n12549), .a(net_9278) );
in01f01  g7062 ( .o(n12550), .a(net_9277) );
in01f01  g7063 ( .o(n12551), .a(net_9276) );
no02f01  g7064 ( .o(n12552), .a(n10001), .b(n10003) );
in01f01  g7065 ( .o(n12553), .a(n12552) );
no02f01  g7066 ( .o(n12554), .a(n12553), .b(n12551) );
in01f01  g7067 ( .o(n12555), .a(n12554) );
no03f01  g7068 ( .o(n12556), .a(n12555), .b(n12550), .c(n12549) );
ao12f01  g7069 ( .o(n12557), .a(net_9278), .b(n12554), .c(net_9277) );
no03f01  g7070 ( .o(n5605), .a(n12557), .b(n12556), .c(n10005) );
in01f01  g7071 ( .o(n12559), .a(_net_10425) );
ao12f01  g7072 ( .o(n12560), .a(n5658), .b(n6052_1), .c(x5143) );
oa12f01  g7073 ( .o(n5610), .a(n12560), .b(n6048), .c(n12559) );
ao12f01  g7074 ( .o(n12562), .a(n5658), .b(n6532), .c(_net_254) );
ao22f01  g7075 ( .o(n12563), .a(n6535), .b(x4520), .c(n6534), .d(net_10014) );
na02f01  g7076 ( .o(n5619), .a(n12563), .b(n12562) );
na02f01  g7077 ( .o(n12565), .a(n6038), .b(net_247) );
na02f01  g7078 ( .o(n12566), .a(n6037_1), .b(net_9876) );
ao22f01  g7079 ( .o(n12567), .a(n6044), .b(x5077), .c(n6042_1), .d(_net_10321) );
na04f01  g7080 ( .o(n5624), .a(n12567), .b(n12566), .c(n12565), .d(n6040) );
ao22f01  g7081 ( .o(n12569), .a(n5842), .b(net_9716), .c(n5841), .d(_net_156) );
na02f01  g7082 ( .o(n12570), .a(n5847), .b(net_10013) );
ao22f01  g7083 ( .o(n12571), .a(n5850), .b(net_9815), .c(n5849_1), .d(net_9914) );
na03f01  g7084 ( .o(n5642), .a(n12571), .b(n12570), .c(n12569) );
ao12f01  g7085 ( .o(n12573), .a(n5658), .b(n6532), .c(net_258) );
ao22f01  g7086 ( .o(n12574), .a(n6535), .b(x4209), .c(n6534), .d(net_10018) );
na02f01  g7087 ( .o(n5647), .a(n12574), .b(n12573) );
no02f01  g7088 ( .o(n12576), .a(n7577), .b(n7582) );
in01f01  g7089 ( .o(n12577), .a(n12576) );
ao12f01  g7090 ( .o(n12578), .a(n12577), .b(n7632), .c(n11572) );
na02f01  g7091 ( .o(n12579), .a(n7632), .b(n11572) );
oa12f01  g7092 ( .o(n12580), .a(n11345), .b(n12576), .c(n12579) );
ao22f01  g7093 ( .o(n12581), .a(n11577), .b(_net_9603), .c(n11576), .d(net_103) );
oa12f01  g7094 ( .o(n5661), .a(n12581), .b(n12580), .c(n12578) );
in01f01  g7095 ( .o(n12583), .a(_net_10212) );
ao12f01  g7096 ( .o(n12584), .a(n5658), .b(n6887), .c(x5364) );
oa12f01  g7097 ( .o(n5666), .a(n12584), .b(n6885_1), .c(n12583) );
ao12f01  g7098 ( .o(n12586), .a(n5658), .b(n5678), .c(net_250) );
ao22f01  g7099 ( .o(n12587), .a(n5681_1), .b(x4851), .c(n5680), .d(net_9713) );
na02f01  g7100 ( .o(n5671), .a(n12587), .b(n12586) );
in01f01  g7101 ( .o(n12589), .a(n10433) );
ao12f01  g7102 ( .o(n12590), .a(n12589), .b(n10430), .c(n8026_1) );
no02f01  g7103 ( .o(n5676), .a(n12590), .b(n7701) );
in01f01  g7104 ( .o(n12592), .a(_net_10094) );
na02f01  g7105 ( .o(n12593), .a(n12592), .b(net_10093) );
ao12f01  g7106 ( .o(n5685), .a(n6155_1), .b(n12593), .c(n10693) );
in01f01  g7107 ( .o(n12595), .a(net_9252) );
oa22f01  g7108 ( .o(n5690), .a(n10323), .b(n12595), .c(n10322), .d(n6089) );
oa22f01  g7109 ( .o(n5695), .a(n5694), .b(n5711), .c(n5692), .d(n5573) );
ao12f01  g7110 ( .o(n12598), .a(n6131_1), .b(n6148), .c(net_9366) );
oa12f01  g7111 ( .o(n5700), .a(n12598), .b(n8101_1), .c(n7104_1) );
na02f01  g7112 ( .o(n12600), .a(n9068), .b(_net_10225) );
na02f01  g7113 ( .o(n5705), .a(n12600), .b(n9070) );
in01f01  g7114 ( .o(n12602), .a(n7039_1) );
no02f01  g7115 ( .o(n12603), .a(n7050), .b(n7008) );
na03f01  g7116 ( .o(n12604), .a(n12603), .b(n7046), .c(n12602) );
in01f01  g7117 ( .o(n12605), .a(n7046) );
in01f01  g7118 ( .o(n12606), .a(n12603) );
oa12f01  g7119 ( .o(n12607), .a(n12606), .b(n12605), .c(n7039_1) );
na02f01  g7120 ( .o(n5710), .a(n12607), .b(n12604) );
na02f01  g7121 ( .o(n12609), .a(net_111), .b(_net_9606) );
na02f01  g7122 ( .o(n12610), .a(n7619), .b(n7561) );
in01f01  g7123 ( .o(n12611), .a(n7621_1) );
na02f01  g7124 ( .o(n12612), .a(n12611), .b(n12610) );
na02f01  g7125 ( .o(n12613), .a(n12612), .b(n7540) );
ao12f01  g7126 ( .o(n12614), .a(n7519_1), .b(n12613), .c(n7523) );
na02f01  g7127 ( .o(n12615), .a(n7514_1), .b(_net_9556) );
in01f01  g7128 ( .o(n12616), .a(n12615) );
no02f01  g7129 ( .o(n12617), .a(n12616), .b(n7522) );
in01f01  g7130 ( .o(n12618), .a(n12617) );
no02f01  g7131 ( .o(n12619), .a(n12618), .b(n12614) );
in01f01  g7132 ( .o(n12620), .a(n7519_1) );
in01f01  g7133 ( .o(n12621), .a(n7540) );
ao12f01  g7134 ( .o(n12622), .a(n12621), .b(n12611), .c(n12610) );
oa12f01  g7135 ( .o(n12623), .a(n12620), .b(n12622), .c(n7524_1) );
oa12f01  g7136 ( .o(n12624), .a(n7500), .b(n12617), .c(n12623) );
oa12f01  g7137 ( .o(n5719), .a(n12609), .b(n12624), .c(n12619) );
no02f01  g7138 ( .o(n12626), .a(n7045), .b(n7013) );
in01f01  g7139 ( .o(n12627), .a(n12626) );
na02f01  g7140 ( .o(n12628), .a(n12627), .b(n7037) );
in01f01  g7141 ( .o(n12629), .a(n7037) );
na02f01  g7142 ( .o(n12630), .a(n12626), .b(n12629) );
na02f01  g7143 ( .o(n5724), .a(n12630), .b(n12628) );
in01f01  g7144 ( .o(n12632), .a(net_10386) );
oa22f01  g7145 ( .o(n5729), .a(n10211), .b(n5597_1), .c(n10210), .d(n12632) );
ao22f01  g7146 ( .o(n12634), .a(n5842), .b(net_9664), .c(n5841), .d(net_102) );
na02f01  g7147 ( .o(n12635), .a(n5847), .b(net_9961) );
ao22f01  g7148 ( .o(n12636), .a(n5850), .b(net_9763), .c(n5849_1), .d(net_9862) );
na03f01  g7149 ( .o(n5734), .a(n12636), .b(n12635), .c(n12634) );
in01f01  g7150 ( .o(n12638), .a(_net_9537) );
no03f01  g7151 ( .o(n12639), .a(n10356), .b(n11533), .c(n12638) );
no04f01  g7152 ( .o(n12640), .a(n12638), .b(_net_9250), .c(_net_9437), .d(n5658) );
na02f01  g7153 ( .o(n12641), .a(_net_9537), .b(n5489) );
oa12f01  g7154 ( .o(n12642), .a(n8399_1), .b(_net_9537), .c(_net_9437) );
oa22f01  g7155 ( .o(n12643), .a(n12642), .b(n5867), .c(n12641), .d(n5871) );
no03f01  g7156 ( .o(n12644), .a(n12643), .b(n12640), .c(n12639) );
no02f01  g7157 ( .o(n12645), .a(n5881), .b(n5876) );
oa12f01  g7158 ( .o(n12646), .a(n12645), .b(n5878_1), .c(_net_9537) );
no02f01  g7159 ( .o(n12647), .a(n12638), .b(_net_9250) );
na02f01  g7160 ( .o(n12648), .a(n12647), .b(n5892) );
na03f01  g7161 ( .o(n5739), .a(n12648), .b(n12646), .c(n12644) );
in01f01  g7162 ( .o(n12650), .a(x3772) );
na02f01  g7163 ( .o(n12651), .a(_net_10278), .b(_net_10277) );
no02f01  g7164 ( .o(n12652), .a(n12651), .b(n11735) );
in01f01  g7165 ( .o(n12653), .a(_net_10279) );
no02f01  g7166 ( .o(n12654), .a(n11736), .b(n12653) );
no03f01  g7167 ( .o(n12655), .a(n12654), .b(n12652), .c(n12650) );
in01f01  g7168 ( .o(n12656), .a(_net_10302) );
ao12f01  g7169 ( .o(n12657), .a(n5658), .b(n12656), .c(_net_10301) );
na02f01  g7170 ( .o(n12658), .a(n12657), .b(x1010) );
oa22f01  g7171 ( .o(n5744), .a(n12658), .b(n12655), .c(n12657), .d(n5658) );
no02f01  g7172 ( .o(n12660), .a(_net_10155), .b(n7771) );
no02f01  g7173 ( .o(n12661), .a(n12660), .b(n7770) );
in01f01  g7174 ( .o(n12662), .a(n12661) );
oa12f01  g7175 ( .o(n12663), .a(n12662), .b(n7789), .c(n7773_1) );
na03f01  g7176 ( .o(n12664), .a(n12661), .b(n7790), .c(n7774) );
na02f01  g7177 ( .o(n5748), .a(n12664), .b(n12663) );
ao12f01  g7178 ( .o(n12666), .a(n7883), .b(n7923), .c(_net_9316) );
oa12f01  g7179 ( .o(n5753), .a(n12666), .b(n7925_1), .c(n8762_1) );
in01f01  g7180 ( .o(n12668), .a(_net_10320) );
ao12f01  g7181 ( .o(n12669), .a(n5658), .b(n5774), .c(x5143) );
oa12f01  g7182 ( .o(n5758), .a(n12669), .b(n5770), .c(n12668) );
na02f01  g7183 ( .o(n12671), .a(n7937), .b(_net_234) );
na02f01  g7184 ( .o(n12672), .a(n7936), .b(net_9764) );
ao22f01  g7185 ( .o(n12673), .a(n7943), .b(_net_10203), .c(n7942), .d(x5901) );
na04f01  g7186 ( .o(n5763), .a(n12673), .b(n12672), .c(n12671), .d(n7939) );
oa22f01  g7187 ( .o(n5768), .a(n5907), .b(n5829), .c(n5905), .d(n5640) );
in01f01  g7188 ( .o(n12676), .a(_net_10419) );
ao12f01  g7189 ( .o(n12677), .a(n5658), .b(n6052_1), .c(x5548) );
oa12f01  g7190 ( .o(n5773), .a(n12677), .b(n6048), .c(n12676) );
in01f01  g7191 ( .o(n12679), .a(net_10285) );
oa22f01  g7192 ( .o(n5782), .a(n9353), .b(n5615), .c(n9352), .d(n12679) );
na02f01  g7193 ( .o(n12681), .a(n6056), .b(net_238) );
na02f01  g7194 ( .o(n12682), .a(n6055), .b(net_9966) );
ao22f01  g7195 ( .o(n12683), .a(n6062_1), .b(x5647), .c(n6060), .d(_net_10417) );
na04f01  g7196 ( .o(n5787), .a(n12683), .b(n12682), .c(n12681), .d(n6058) );
na03f01  g7197 ( .o(n12685), .a(n8748), .b(n7974), .c(_net_9638) );
no02f01  g7198 ( .o(n12686), .a(n7969), .b(n7964) );
ao12f01  g7199 ( .o(n12687), .a(n8751), .b(n12686), .c(n12685) );
na03f01  g7200 ( .o(n12688), .a(n9542), .b(_net_9638), .c(_net_9641) );
na02f01  g7201 ( .o(n12689), .a(n9495), .b(_net_9638) );
no04f01  g7202 ( .o(n12690), .a(n8773), .b(net_9612), .c(n8784), .d(n8772_1) );
ao12f01  g7203 ( .o(n12691), .a(n12690), .b(n9496), .c(_net_9638) );
na03f01  g7204 ( .o(n12692), .a(n12691), .b(n12689), .c(n12688) );
no02f01  g7205 ( .o(n12693), .a(n12692), .b(n12687) );
no02f01  g7206 ( .o(n5792), .a(n12693), .b(n9500) );
na02f01  g7207 ( .o(n12695), .a(n6038), .b(net_248) );
na02f01  g7208 ( .o(n12696), .a(n6037_1), .b(net_9877) );
ao22f01  g7209 ( .o(n12697), .a(n6044), .b(x5003), .c(n6042_1), .d(_net_10322) );
na04f01  g7210 ( .o(n5797), .a(n12697), .b(n12696), .c(n12695), .d(n6040) );
oa22f01  g7211 ( .o(n5802), .a(n5907), .b(n8605), .c(n5905), .d(n5597_1) );
in01f01  g7212 ( .o(n12700), .a(n7908) );
ao12f01  g7213 ( .o(n12701), .a(n9767), .b(n9756), .c(n7732) );
ao12f01  g7214 ( .o(n12702), .a(n9759), .b(n12701), .c(n12700) );
no02f01  g7215 ( .o(n12703), .a(n9767), .b(n7732) );
oa12f01  g7216 ( .o(n12704), .a(_net_9355), .b(n8754), .c(net_9151) );
no02f01  g7217 ( .o(n12705), .a(n7734_1), .b(n9767) );
ao22f01  g7218 ( .o(n12706), .a(n12705), .b(n9772), .c(n9774), .d(_net_9355) );
oa12f01  g7219 ( .o(n12707), .a(n12706), .b(n12704), .c(n9769) );
ao12f01  g7220 ( .o(n12708), .a(n12707), .b(n12703), .c(n9766) );
oa12f01  g7221 ( .o(n5807), .a(n12708), .b(n12702), .c(n9760) );
na03f01  g7222 ( .o(n12710), .a(n9061), .b(n8969), .c(n8957) );
na04f01  g7223 ( .o(n12711), .a(n9172), .b(n9220), .c(n9180), .d(n8978) );
no04f01  g7224 ( .o(n12712), .a(n12711), .b(n12710), .c(_net_10225), .d(_net_10226) );
no03f01  g7225 ( .o(n5820), .a(n12712), .b(_net_9851), .c(n9385) );
na02f01  g7226 ( .o(n12714), .a(n8200_1), .b(n9129) );
no02f01  g7227 ( .o(n12715), .a(_net_9926), .b(n9129) );
oa12f01  g7228 ( .o(n12716), .a(n8183), .b(n12715), .c(n9095) );
na02f01  g7229 ( .o(n12717), .a(n8202), .b(_net_10350) );
na03f01  g7230 ( .o(n5825), .a(n12717), .b(n12716), .c(n12714) );
na02f01  g7231 ( .o(n12719), .a(n5577), .b(n7991) );
in01f01  g7232 ( .o(n12720), .a(n9461) );
no02f01  g7233 ( .o(n12721), .a(n9460), .b(n9459) );
oa12f01  g7234 ( .o(n12722), .a(n7998), .b(n12721), .c(n12720) );
no02f01  g7235 ( .o(n12723), .a(n8002), .b(n9459) );
no02f01  g7236 ( .o(n12724), .a(n12723), .b(n5658) );
na03f01  g7237 ( .o(n5830), .a(n12724), .b(n12722), .c(n12719) );
in01f01  g7238 ( .o(n12726), .a(n8047) );
oa22f01  g7239 ( .o(n12727), .a(n12726), .b(n10462), .c(n6563), .d(n10818) );
ao12f01  g7240 ( .o(n12728), .a(n12727), .b(n6555), .c(net_9984) );
ao22f01  g7241 ( .o(n12729), .a(n6573), .b(net_9885), .c(n6572), .d(net_10387) );
ao22f01  g7242 ( .o(n12730), .a(n6602), .b(net_10016), .c(n6577), .d(net_9687) );
na02f01  g7243 ( .o(n12731), .a(n6584_1), .b(net_9786) );
ao22f01  g7244 ( .o(n12732), .a(n6599_1), .b(net_9849), .c(n6582), .d(net_9917) );
na02f01  g7245 ( .o(n12733), .a(n12732), .b(n12731) );
ao22f01  g7246 ( .o(n12734), .a(n6592), .b(net_10177), .c(n6590), .d(net_10047) );
ao22f01  g7247 ( .o(n12735), .a(n6597), .b(net_9750), .c(n6585), .d(net_9719) );
ao22f01  g7248 ( .o(n12736), .a(n6603), .b(net_10492), .c(n6580), .d(net_9818) );
ao22f01  g7249 ( .o(n12737), .a(n6606), .b(net_9948), .c(n6605), .d(net_10282) );
na04f01  g7250 ( .o(n12738), .a(n12737), .b(n12736), .c(n12735), .d(n12734) );
no02f01  g7251 ( .o(n12739), .a(n12738), .b(n12733) );
na04f01  g7252 ( .o(n5835), .a(n12739), .b(n12730), .c(n12729), .d(n12728) );
na02f01  g7253 ( .o(n12741), .a(n6038), .b(net_239) );
na02f01  g7254 ( .o(n12742), .a(n6037_1), .b(net_9868) );
ao22f01  g7255 ( .o(n12743), .a(n6044), .b(x5601), .c(n6042_1), .d(_net_10313) );
na04f01  g7256 ( .o(n5839), .a(n12743), .b(n12742), .c(n12741), .d(n6040) );
oa22f01  g7257 ( .o(n5844), .a(n7738_1), .b(n6457), .c(n7736), .d(n8984) );
ao22f01  g7258 ( .o(n12746), .a(n5702), .b(x2707), .c(n5701), .d(_net_9398) );
oa12f01  g7259 ( .o(n5849), .a(n12746), .b(n5700_1), .c(n5737) );
ao12f01  g7260 ( .o(n12748), .a(n8890), .b(n8881), .c(n8856) );
no02f01  g7261 ( .o(n12749), .a(n12748), .b(n8907) );
no02f01  g7262 ( .o(n12750), .a(n8899), .b(n8884) );
na02f01  g7263 ( .o(n12751), .a(n12750), .b(n12749) );
in01f01  g7264 ( .o(n12752), .a(n12750) );
oa12f01  g7265 ( .o(n12753), .a(n12752), .b(n12748), .c(n8907) );
na02f01  g7266 ( .o(n5858), .a(n12753), .b(n12751) );
na02f01  g7267 ( .o(n12755), .a(n6038), .b(net_258) );
na02f01  g7268 ( .o(n12756), .a(n6037_1), .b(net_9887) );
ao22f01  g7269 ( .o(n12757), .a(n6044), .b(x4209), .c(n6042_1), .d(_net_10332) );
na04f01  g7270 ( .o(n5863), .a(n12757), .b(n12756), .c(n12755), .d(n6040) );
in01f01  g7271 ( .o(n12759), .a(_net_9187) );
oa22f01  g7272 ( .o(n5868), .a(n8349_1), .b(n8017), .c(n8347), .d(n12759) );
no02f01  g7273 ( .o(n12761), .a(n5751), .b(_net_10118) );
in01f01  g7274 ( .o(n12762), .a(n12761) );
na02f01  g7275 ( .o(n12763), .a(n5751), .b(_net_10118) );
na02f01  g7276 ( .o(n5873), .a(n12763), .b(n12762) );
ao12f01  g7277 ( .o(n12765), .a(n5658), .b(n6887), .c(x4694) );
oa12f01  g7278 ( .o(n5878), .a(n12765), .b(n6885_1), .c(n8957) );
ao12f01  g7279 ( .o(n12767), .a(n5658), .b(n5678), .c(net_244) );
ao22f01  g7280 ( .o(n12768), .a(n5681_1), .b(x5289), .c(n5680), .d(net_9707) );
na02f01  g7281 ( .o(n5883), .a(n12768), .b(n12767) );
in01f01  g7282 ( .o(n12770), .a(_net_10412) );
ao12f01  g7283 ( .o(n12771), .a(n5658), .b(n6052_1), .c(x5961) );
oa12f01  g7284 ( .o(n5888), .a(n12771), .b(n6048), .c(n12770) );
na02f01  g7285 ( .o(n12773), .a(n6056), .b(net_252) );
na02f01  g7286 ( .o(n12774), .a(n6055), .b(net_9980) );
ao22f01  g7287 ( .o(n12775), .a(n6062_1), .b(x4694), .c(n6060), .d(_net_10431) );
na04f01  g7288 ( .o(n5893), .a(n12775), .b(n12774), .c(n12773), .d(n6058) );
in01f01  g7289 ( .o(n12777), .a(_net_10097) );
ao12f01  g7290 ( .o(n12778), .a(n5658), .b(n6160_1), .c(x5961) );
oa12f01  g7291 ( .o(n5898), .a(n12778), .b(n6159), .c(n12777) );
na02f01  g7292 ( .o(n12780), .a(net_10404), .b(net_10390) );
ao22f01  g7293 ( .o(n12781), .a(net_10391), .b(net_10405), .c(net_10389), .d(net_10403) );
ao22f01  g7294 ( .o(n12782), .a(net_10389), .b(net_10402), .c(net_10399), .d(net_10386) );
ao22f01  g7295 ( .o(n12783), .a(net_10388), .b(net_10401), .c(net_10400), .d(net_10387) );
na04f01  g7296 ( .o(n5903), .a(n12783), .b(n12782), .c(n12781), .d(n12780) );
in01f01  g7297 ( .o(n12785), .a(_net_10102) );
ao12f01  g7298 ( .o(n12786), .a(n5658), .b(n6160_1), .c(x5647) );
oa12f01  g7299 ( .o(n5908), .a(n12786), .b(n6159), .c(n12785) );
no02f01  g7300 ( .o(n12788), .a(n6919_1), .b(n6910_1) );
in01f01  g7301 ( .o(n12789), .a(n12788) );
ao12f01  g7302 ( .o(n12790), .a(n6933), .b(n12789), .c(n6909) );
oa12f01  g7303 ( .o(n12791), .a(n12790), .b(n12789), .c(n6909) );
na02f01  g7304 ( .o(n12792), .a(n6938), .b(_net_10261) );
na02f01  g7305 ( .o(n12793), .a(n12792), .b(n6940) );
ao22f01  g7306 ( .o(n12794), .a(n12793), .b(n6175), .c(n6168), .d(_net_10261) );
na02f01  g7307 ( .o(n5913), .a(n12794), .b(n12791) );
oa22f01  g7308 ( .o(n5921), .a(n6989_1), .b(n5612), .c(n6988), .d(n9238) );
na02f01  g7309 ( .o(n12797), .a(n7937), .b(net_253) );
na02f01  g7310 ( .o(n12798), .a(n7936), .b(net_9783) );
ao22f01  g7311 ( .o(n12799), .a(n7943), .b(_net_10222), .c(n7942), .d(x4587) );
na04f01  g7312 ( .o(n5926), .a(n12799), .b(n12798), .c(n12797), .d(n7939) );
no02f01  g7313 ( .o(n12801), .a(n6903), .b(n6785) );
no02f01  g7314 ( .o(n12802), .a(n6908), .b(n12801) );
no02f01  g7315 ( .o(n12803), .a(_net_9830), .b(_net_10260) );
no02f01  g7316 ( .o(n12804), .a(n6904), .b(n6902) );
no02f01  g7317 ( .o(n12805), .a(n12804), .b(n12803) );
in01f01  g7318 ( .o(n12806), .a(n12805) );
ao12f01  g7319 ( .o(n12807), .a(n6933), .b(n12806), .c(n12802) );
oa12f01  g7320 ( .o(n12808), .a(n12807), .b(n12806), .c(n12802) );
oa12f01  g7321 ( .o(n12809), .a(_net_10260), .b(n6936), .c(_net_10259) );
ao12f01  g7322 ( .o(n12810), .a(n6846_1), .b(n12809), .c(n6938) );
ao12f01  g7323 ( .o(n12811), .a(n12810), .b(n6168), .c(_net_10260) );
na02f01  g7324 ( .o(n5931), .a(n12811), .b(n12808) );
oa22f01  g7325 ( .o(n5944), .a(n8418), .b(n8736), .c(n8417), .d(n5561) );
ao12f01  g7326 ( .o(n12814), .a(n5658), .b(n5678), .c(net_248) );
ao22f01  g7327 ( .o(n12815), .a(n5681_1), .b(x5003), .c(n5680), .d(net_9711) );
na02f01  g7328 ( .o(n5949), .a(n12815), .b(n12814) );
in01f01  g7329 ( .o(n12817), .a(net_9726) );
oa22f01  g7330 ( .o(n5954), .a(n7367), .b(n12817), .c(n7365_1), .d(n5570) );
na02f01  g7331 ( .o(n12819), .a(n8234), .b(n8221) );
no02f01  g7332 ( .o(n12820), .a(n8219_1), .b(_net_10470) );
no02f01  g7333 ( .o(n12821), .a(n12820), .b(n8218) );
in01f01  g7334 ( .o(n12822), .a(n12821) );
na02f01  g7335 ( .o(n12823), .a(n12822), .b(n12819) );
na03f01  g7336 ( .o(n12824), .a(n12821), .b(n8234), .c(n8221) );
na02f01  g7337 ( .o(n5959), .a(n12824), .b(n12823) );
ao12f01  g7338 ( .o(n12826), .a(n5658), .b(n7844), .c(net_244) );
ao22f01  g7339 ( .o(n12827), .a(n7847), .b(x5289), .c(n7846), .d(net_9806) );
na02f01  g7340 ( .o(n5964), .a(n12827), .b(n12826) );
no02f01  g7341 ( .o(n12829), .a(n7524_1), .b(n7519_1) );
in01f01  g7342 ( .o(n12830), .a(n12829) );
na02f01  g7343 ( .o(n12831), .a(n12830), .b(n12613) );
na02f01  g7344 ( .o(n12832), .a(n12829), .b(n12622) );
na02f01  g7345 ( .o(n5969), .a(n12832), .b(n12831) );
oa22f01  g7346 ( .o(n5978), .a(n7756), .b(n6367), .c(n7755), .d(n12253) );
oa22f01  g7347 ( .o(n12835), .a(n8841), .b(n7593), .c(n6024), .d(n6025) );
na02f01  g7348 ( .o(n12836), .a(n6024), .b(n6025) );
oa22f01  g7349 ( .o(n12837), .a(n7072), .b(n7073_1), .c(n6625), .d(n7571_1) );
ao12f01  g7350 ( .o(n12838), .a(n12837), .b(n12836), .c(n12835) );
oa12f01  g7351 ( .o(n12839), .a(n7571_1), .b(n7072), .c(n7073_1) );
oa22f01  g7352 ( .o(n12840), .a(n12839), .b(n5938), .c(n5941), .d(_net_9293) );
oa22f01  g7353 ( .o(n12841), .a(n6634_1), .b(n7545), .c(n6614_1), .d(n7552_1) );
oa22f01  g7354 ( .o(n12842), .a(n5976), .b(n8469), .c(n6617), .d(n7605_1) );
no02f01  g7355 ( .o(n12843), .a(n12842), .b(n12841) );
oa12f01  g7356 ( .o(n12844), .a(n12843), .b(n12840), .c(n12838) );
oa12f01  g7357 ( .o(n12845), .a(n7605_1), .b(n5976), .c(n8469) );
no03f01  g7358 ( .o(n12846), .a(n12845), .b(n12841), .c(n5965) );
no03f01  g7359 ( .o(n12847), .a(n12841), .b(n5968), .c(_net_9295) );
oa12f01  g7360 ( .o(n12848), .a(n7545), .b(n6614_1), .c(n7552_1) );
oa22f01  g7361 ( .o(n12849), .a(n12848), .b(n5961), .c(n5958), .d(_net_9297) );
no03f01  g7362 ( .o(n12850), .a(n12849), .b(n12847), .c(n12846) );
ao22f01  g7363 ( .o(n12851), .a(n5997), .b(_net_9298), .c(n5993_1), .d(_net_9299) );
na02f01  g7364 ( .o(n12852), .a(n5986), .b(_net_9300) );
na02f01  g7365 ( .o(n12853), .a(n12852), .b(n12851) );
ao12f01  g7366 ( .o(n12854), .a(n12853), .b(n12850), .c(n12844) );
no02f01  g7367 ( .o(n12855), .a(n5994), .b(n7529_1) );
no03f01  g7368 ( .o(n12856), .a(n12855), .b(n5997), .c(_net_9298) );
oa22f01  g7369 ( .o(n12857), .a(n5993_1), .b(_net_9299), .c(n5986), .d(_net_9300) );
oa12f01  g7370 ( .o(n12858), .a(n12852), .b(n12857), .c(n12856) );
no02f01  g7371 ( .o(n12859), .a(n6017), .b(n6011) );
na04f01  g7372 ( .o(n12860), .a(n12859), .b(n12858), .c(n8918), .d(net_9288) );
no02f01  g7373 ( .o(n5983), .a(n12860), .b(n12854) );
in01f01  g7374 ( .o(n12862), .a(net_10509) );
na02f01  g7375 ( .o(n12863), .a(net_263), .b(net_10490) );
ao12f01  g7376 ( .o(n5988), .a(n9667), .b(n12863), .c(n12862) );
na02f01  g7377 ( .o(n12865), .a(n7937), .b(net_242) );
na02f01  g7378 ( .o(n12866), .a(n7936), .b(net_9772) );
ao22f01  g7379 ( .o(n12867), .a(n7943), .b(_net_10211), .c(n7942), .d(x5427) );
na04f01  g7380 ( .o(n5993), .a(n12867), .b(n12866), .c(n12865), .d(n7939) );
na02f01  g7381 ( .o(n12869), .a(n6349), .b(n6345) );
na02f01  g7382 ( .o(n12870), .a(n6351_1), .b(_net_9267) );
oa12f01  g7383 ( .o(n6005), .a(n12870), .b(n12869), .c(n6348) );
in01f01  g7384 ( .o(n12872), .a(n9215) );
no02f01  g7385 ( .o(n12873), .a(n9176), .b(n9173) );
na03f01  g7386 ( .o(n12874), .a(n12873), .b(n12872), .c(n9178) );
in01f01  g7387 ( .o(n12875), .a(n12873) );
oa12f01  g7388 ( .o(n12876), .a(n12875), .b(n9215), .c(n9177) );
na02f01  g7389 ( .o(n6013), .a(n12876), .b(n12874) );
na02f01  g7390 ( .o(n12878), .a(n6750), .b(n6751) );
no02f01  g7391 ( .o(n12879), .a(n6751), .b(_net_9728) );
oa12f01  g7392 ( .o(n12880), .a(n10948), .b(n12879), .c(n6728_1) );
na02f01  g7393 ( .o(n12881), .a(n6760), .b(_net_10140) );
na03f01  g7394 ( .o(n6018), .a(n12881), .b(n12880), .c(n12878) );
na02f01  g7395 ( .o(n12883), .a(net_10500), .b(net_10507) );
ao22f01  g7396 ( .o(n12884), .a(net_10505), .b(net_10498), .c(net_10499), .d(net_10506) );
ao22f01  g7397 ( .o(n12885), .a(net_10500), .b(net_10508), .c(net_10509), .d(net_10501) );
ao22f01  g7398 ( .o(n12886), .a(net_10504), .b(net_10497), .c(net_10510), .d(net_10502) );
na04f01  g7399 ( .o(n6023), .a(n12886), .b(n12885), .c(n12884), .d(n12883) );
na02f01  g7400 ( .o(n12888), .a(n7358), .b(net_258) );
na02f01  g7401 ( .o(n12889), .a(n7352), .b(net_9689) );
ao22f01  g7402 ( .o(n12890), .a(n7357), .b(_net_10122), .c(n7353), .d(x4209) );
na04f01  g7403 ( .o(n6028), .a(n12890), .b(n12889), .c(n12888), .d(n7355_1) );
na02f01  g7404 ( .o(n12892), .a(n10775), .b(n6697) );
oa22f01  g7405 ( .o(n6037), .a(n12892), .b(n6688), .c(n6685), .d(n6691) );
no03f01  g7406 ( .o(n12894), .a(n10304), .b(n10303), .c(n9720) );
in01f01  g7407 ( .o(n12895), .a(n12894) );
no02f01  g7408 ( .o(n12896), .a(n10305), .b(n10302) );
ao12f01  g7409 ( .o(n12897), .a(n7875), .b(n12896), .c(n12895) );
oa12f01  g7410 ( .o(n12898), .a(n12897), .b(n12896), .c(n12895) );
na02f01  g7411 ( .o(n12899), .a(n9733), .b(n9037) );
no02f01  g7412 ( .o(n12900), .a(n11333), .b(n7451_1) );
ao22f01  g7413 ( .o(n12901), .a(n12900), .b(n12899), .c(n7453), .d(_net_10462) );
na02f01  g7414 ( .o(n6042), .a(n12901), .b(n12898) );
na02f01  g7415 ( .o(n12903), .a(n1792), .b(n7991) );
na02f01  g7416 ( .o(n12904), .a(n9465), .b(net_9526) );
ao12f01  g7417 ( .o(n12905), .a(n7999), .b(n12904), .c(n9567) );
in01f01  g7418 ( .o(n12906), .a(net_9526) );
oa12f01  g7419 ( .o(n12907), .a(x6599), .b(n8002), .c(n12906) );
no02f01  g7420 ( .o(n12908), .a(n12907), .b(n12905) );
na02f01  g7421 ( .o(n6047), .a(n12908), .b(n12903) );
no02f01  g7422 ( .o(n12910), .a(n8265), .b(_net_201) );
na02f01  g7423 ( .o(n12911), .a(n8268_1), .b(n573) );
oa22f01  g7424 ( .o(n6052), .a(n12911), .b(n12910), .c(n8280), .d(n8259) );
ao22f01  g7425 ( .o(n12913), .a(n5842), .b(net_9720), .c(n5841), .d(_net_160) );
na02f01  g7426 ( .o(n12914), .a(n5847), .b(net_10017) );
ao22f01  g7427 ( .o(n12915), .a(n5850), .b(net_9819), .c(n5849_1), .d(net_9918) );
na03f01  g7428 ( .o(n6057), .a(n12915), .b(n12914), .c(n12913) );
oa22f01  g7429 ( .o(n6062), .a(n7480_1), .b(n6799), .c(n7478), .d(n5606) );
ao22f01  g7430 ( .o(n12918), .a(n5842), .b(_net_9735), .c(n5841), .d(_net_176) );
na02f01  g7431 ( .o(n12919), .a(n5847), .b(_net_10032) );
ao22f01  g7432 ( .o(n12920), .a(n5850), .b(_net_9834), .c(n5849_1), .d(_net_9933) );
na03f01  g7433 ( .o(n6072), .a(n12920), .b(n12919), .c(n12918) );
in01f01  g7434 ( .o(n12922), .a(net_10510) );
na02f01  g7435 ( .o(n12923), .a(_net_9117), .b(net_10490) );
ao12f01  g7436 ( .o(n6077), .a(n9667), .b(n12923), .c(n12922) );
na02f01  g7437 ( .o(n12925), .a(n6038), .b(net_237) );
na02f01  g7438 ( .o(n12926), .a(n6037_1), .b(net_9866) );
ao22f01  g7439 ( .o(n12927), .a(n6044), .b(x5722), .c(n6042_1), .d(_net_10311) );
na04f01  g7440 ( .o(n6082), .a(n12927), .b(n12926), .c(n12925), .d(n6040) );
ao22f01  g7441 ( .o(n12929), .a(n5842), .b(net_9707), .c(n5841), .d(net_147) );
na02f01  g7442 ( .o(n12930), .a(n5847), .b(net_10004) );
ao22f01  g7443 ( .o(n12931), .a(n5850), .b(net_9806), .c(n5849_1), .d(net_9905) );
na03f01  g7444 ( .o(n6087), .a(n12931), .b(n12930), .c(n12929) );
ao22f01  g7445 ( .o(n12933), .a(n6602), .b(net_10003), .c(n6597), .d(net_9738) );
ao22f01  g7446 ( .o(n12934), .a(n6577), .b(net_9674), .c(n6555), .d(net_9971) );
in01f01  g7447 ( .o(n12935), .a(net_9805) );
oa22f01  g7448 ( .o(n12936), .a(n6966_1), .b(n11884), .c(n9978), .d(n12935) );
na02f01  g7449 ( .o(n12937), .a(n6585), .b(net_9706) );
na02f01  g7450 ( .o(n12938), .a(n6582), .b(net_9904) );
na02f01  g7451 ( .o(n12939), .a(n12938), .b(n12937) );
ao22f01  g7452 ( .o(n12940), .a(n6590), .b(net_10035), .c(n6573), .d(net_9872) );
ao22f01  g7453 ( .o(n12941), .a(n6599_1), .b(net_9837), .c(n6584_1), .d(net_9773) );
na02f01  g7454 ( .o(n12942), .a(n12941), .b(n12940) );
no03f01  g7455 ( .o(n12943), .a(n12942), .b(n12939), .c(n12936) );
na03f01  g7456 ( .o(n6107), .a(n12943), .b(n12934), .c(n12933) );
ao12f01  g7457 ( .o(n12945), .a(n5658), .b(n5678), .c(net_258) );
ao22f01  g7458 ( .o(n12946), .a(n5681_1), .b(x4209), .c(n5680), .d(net_9721) );
na02f01  g7459 ( .o(n6111), .a(n12946), .b(n12945) );
in01f01  g7460 ( .o(n12948), .a(_net_10424) );
ao12f01  g7461 ( .o(n12949), .a(n5658), .b(n6052_1), .c(x5225) );
oa12f01  g7462 ( .o(n6116), .a(n12949), .b(n6048), .c(n12948) );
na02f01  g7463 ( .o(n12951), .a(n8939), .b(_net_10330) );
na02f01  g7464 ( .o(n6121), .a(n12951), .b(n8941) );
na02f01  g7465 ( .o(n12953), .a(n7937), .b(_net_254) );
na02f01  g7466 ( .o(n12954), .a(n7936), .b(net_9784) );
ao22f01  g7467 ( .o(n12955), .a(n7943), .b(_net_10223), .c(n7942), .d(x4520) );
na04f01  g7468 ( .o(n6126), .a(n12955), .b(n12954), .c(n12953), .d(n7939) );
na02f01  g7469 ( .o(n12957), .a(n8868), .b(n8846) );
no02f01  g7470 ( .o(n12958), .a(n8871), .b(n8867_1) );
in01f01  g7471 ( .o(n12959), .a(n12958) );
na02f01  g7472 ( .o(n12960), .a(n12959), .b(n12957) );
na03f01  g7473 ( .o(n12961), .a(n12958), .b(n8868), .c(n8846) );
na02f01  g7474 ( .o(n6131), .a(n12961), .b(n12960) );
na02f01  g7475 ( .o(n12963), .a(n8945), .b(_net_10333) );
na02f01  g7476 ( .o(n6141), .a(n12963), .b(n8947) );
na02f01  g7477 ( .o(n12965), .a(n7453), .b(_net_10456) );
na02f01  g7478 ( .o(n12966), .a(n9014), .b(n9013) );
na03f01  g7479 ( .o(n12967), .a(n12966), .b(n9727), .c(n7450) );
in01f01  g7480 ( .o(n12968), .a(n9709) );
in01f01  g7481 ( .o(n12969), .a(n9710) );
na03f01  g7482 ( .o(n12970), .a(n12969), .b(n12968), .c(n9708) );
in01f01  g7483 ( .o(n12971), .a(n9708) );
oa12f01  g7484 ( .o(n12972), .a(n9709), .b(n9710), .c(n12971) );
na03f01  g7485 ( .o(n12973), .a(n12972), .b(n12970), .c(n7431) );
na03f01  g7486 ( .o(n6150), .a(n12973), .b(n12967), .c(n12965) );
no02f01  g7487 ( .o(n12975), .a(n8175_1), .b(n8158) );
no02f01  g7488 ( .o(n12976), .a(n8155_1), .b(n8157) );
in01f01  g7489 ( .o(n12977), .a(n12976) );
ao12f01  g7490 ( .o(n12978), .a(n8184), .b(n12977), .c(n12975) );
oa12f01  g7491 ( .o(n12979), .a(n12978), .b(n12977), .c(n12975) );
na02f01  g7492 ( .o(n12980), .a(n8192), .b(_net_10367) );
na02f01  g7493 ( .o(n12981), .a(n12980), .b(n8194) );
ao22f01  g7494 ( .o(n12982), .a(n12981), .b(n8200_1), .c(n8202), .d(_net_10367) );
na02f01  g7495 ( .o(n6155), .a(n12982), .b(n12979) );
ao22f01  g7496 ( .o(n12984), .a(n5842), .b(net_9699), .c(n5841), .d(net_139) );
na02f01  g7497 ( .o(n12985), .a(n5847), .b(net_9996) );
ao22f01  g7498 ( .o(n12986), .a(n5850), .b(net_9798), .c(n5849_1), .d(net_9897) );
na03f01  g7499 ( .o(n6160), .a(n12986), .b(n12985), .c(n12984) );
ao22f01  g7500 ( .o(n12988), .a(n5842), .b(net_9753), .c(n5841), .d(_net_189) );
na02f01  g7501 ( .o(n12989), .a(n5847), .b(net_10050) );
ao22f01  g7502 ( .o(n12990), .a(n5850), .b(net_9852), .c(n5849_1), .d(net_9951) );
na03f01  g7503 ( .o(n6164), .a(n12990), .b(n12989), .c(n12988) );
oa22f01  g7504 ( .o(n6173), .a(n7367), .b(n9655), .c(n7365_1), .d(n5637) );
na02f01  g7505 ( .o(n12993), .a(n7666), .b(_net_10432) );
na02f01  g7506 ( .o(n6186), .a(n12993), .b(n7668) );
oa22f01  g7507 ( .o(n6191), .a(n7367), .b(n8532), .c(n7365_1), .d(n5606) );
in01f01  g7508 ( .o(n12996), .a(net_10191) );
na02f01  g7509 ( .o(n12997), .a(net_10175), .b(net_264) );
ao12f01  g7510 ( .o(n6196), .a(n8577_1), .b(n12997), .c(n12996) );
na02f01  g7511 ( .o(n12999), .a(n5757), .b(_net_10122) );
na02f01  g7512 ( .o(n6201), .a(n12999), .b(n5759) );
oa22f01  g7513 ( .o(n6206), .a(n5694), .b(n5705_1), .c(n5692), .d(n5585_1) );
na02f01  g7514 ( .o(n13002), .a(n6056), .b(net_249) );
na02f01  g7515 ( .o(n13003), .a(n6055), .b(net_9977) );
ao22f01  g7516 ( .o(n13004), .a(n6062_1), .b(x4937), .c(n6060), .d(_net_10428) );
na04f01  g7517 ( .o(n6211), .a(n13004), .b(n13003), .c(n13002), .d(n6058) );
no02f01  g7518 ( .o(n13006), .a(n9820), .b(_net_9299) );
na02f01  g7519 ( .o(n13007), .a(n9821), .b(n8809_1) );
oa22f01  g7520 ( .o(n6216), .a(n13007), .b(n13006), .c(n8817), .d(n7529_1) );
oa22f01  g7521 ( .o(n6221), .a(n5907), .b(n7429), .c(n5905), .d(n5582_1) );
oa22f01  g7522 ( .o(n6226), .a(n7480_1), .b(n9826), .c(n7478), .d(n5603) );
in01f01  g7523 ( .o(n13011), .a(n7800) );
no03f01  g7524 ( .o(n13012), .a(n7809), .b(n7806_1), .c(n13011) );
in01f01  g7525 ( .o(n13013), .a(n13012) );
no02f01  g7526 ( .o(n13014), .a(n7810), .b(n7766) );
in01f01  g7527 ( .o(n13015), .a(n13014) );
na02f01  g7528 ( .o(n13016), .a(n13015), .b(n13013) );
na02f01  g7529 ( .o(n13017), .a(n13014), .b(n13012) );
na02f01  g7530 ( .o(n6231), .a(n13017), .b(n13016) );
na02f01  g7531 ( .o(n13019), .a(n7453), .b(_net_10457) );
na02f01  g7532 ( .o(n13020), .a(n9727), .b(n9018) );
na03f01  g7533 ( .o(n13021), .a(n13020), .b(n9729), .c(n7450) );
no02f01  g7534 ( .o(n13022), .a(n9707), .b(n9704) );
in01f01  g7535 ( .o(n13023), .a(n13022) );
na02f01  g7536 ( .o(n13024), .a(n13023), .b(n9712) );
na02f01  g7537 ( .o(n13025), .a(n13022), .b(n9711) );
na03f01  g7538 ( .o(n13026), .a(n13025), .b(n13024), .c(n7431) );
na03f01  g7539 ( .o(n6244), .a(n13026), .b(n13021), .c(n13019) );
in01f01  g7540 ( .o(n13028), .a(net_10044) );
no02f01  g7541 ( .o(n13029), .a(n8624), .b(n5658) );
oa12f01  g7542 ( .o(n13030), .a(n13029), .b(n5906), .c(x4587) );
oa12f01  g7543 ( .o(n6249), .a(n13030), .b(n8625), .c(n13028) );
ao12f01  g7544 ( .o(n13032), .a(n5658), .b(n5678), .c(net_236) );
ao22f01  g7545 ( .o(n13033), .a(n5681_1), .b(x5790), .c(n5680), .d(net_9699) );
na02f01  g7546 ( .o(n6258), .a(n13033), .b(n13032) );
in01f01  g7547 ( .o(n13035), .a(_net_10416) );
ao12f01  g7548 ( .o(n13036), .a(n5658), .b(n6052_1), .c(x5722) );
oa12f01  g7549 ( .o(n6263), .a(n13036), .b(n6048), .c(n13035) );
oa22f01  g7550 ( .o(n6268), .a(n5907), .b(n7396), .c(n5905), .d(n5540) );
in01f01  g7551 ( .o(n13039), .a(_net_10321) );
ao12f01  g7552 ( .o(n13040), .a(n5658), .b(n5774), .c(x5077) );
oa12f01  g7553 ( .o(n6277), .a(n13040), .b(n5770), .c(n13039) );
oa22f01  g7554 ( .o(n6282), .a(n5694), .b(n5812_1), .c(n5692), .d(n5552_1) );
na02f01  g7555 ( .o(n13043), .a(_net_10430), .b(n1032) );
na02f01  g7556 ( .o(n13044), .a(n8227_1), .b(_net_10429) );
na02f01  g7557 ( .o(n6287), .a(n13044), .b(n13043) );
ao12f01  g7558 ( .o(n13046), .a(n5658), .b(n6532), .c(_net_231) );
ao22f01  g7559 ( .o(n13047), .a(n6535), .b(x6102), .c(n6534), .d(net_9991) );
na02f01  g7560 ( .o(n6292), .a(n13047), .b(n13046) );
na03f01  g7561 ( .o(n13049), .a(n5880), .b(n5879), .c(net_9535) );
in01f01  g7562 ( .o(n13050), .a(net_9535) );
no03f01  g7563 ( .o(n13051), .a(n8404_1), .b(n13050), .c(_net_9503) );
ao12f01  g7564 ( .o(n13052), .a(net_9544), .b(net_9535), .c(n5883_1) );
no03f01  g7565 ( .o(n13053), .a(n13052), .b(n5886), .c(_net_9250) );
no03f01  g7566 ( .o(n13054), .a(n13050), .b(_net_9437), .c(n5658) );
no03f01  g7567 ( .o(n13055), .a(n13054), .b(n13053), .c(n13051) );
no03f01  g7568 ( .o(n13056), .a(n13050), .b(_net_9250), .c(_net_9437) );
no02f01  g7569 ( .o(n13057), .a(n10356), .b(n13050) );
ao22f01  g7570 ( .o(n13058), .a(n13057), .b(n5857), .c(n13056), .d(n8412) );
na03f01  g7571 ( .o(n6297), .a(n13058), .b(n13055), .c(n13049) );
na03f01  g7572 ( .o(n13060), .a(n6860), .b(_net_9239), .c(_net_9236) );
na02f01  g7573 ( .o(n13061), .a(n6471), .b(_net_9239) );
oa12f01  g7574 ( .o(n13062), .a(n13060), .b(n13061), .c(n7862_1) );
ao12f01  g7575 ( .o(n13063), .a(n13061), .b(n7863), .c(n7852) );
no02f01  g7576 ( .o(n13064), .a(n13063), .b(n13062) );
no03f01  g7577 ( .o(n13065), .a(n7482), .b(n6485), .c(n6491) );
ao12f01  g7578 ( .o(n13066), .a(n6468), .b(n6464_1), .c(_net_9239) );
no03f01  g7579 ( .o(n13067), .a(n13066), .b(n6472), .c(n6463) );
ao22f01  g7580 ( .o(n13068), .a(n10426), .b(n6677), .c(n6476), .d(_net_9239) );
na02f01  g7581 ( .o(n13069), .a(n6491), .b(n8508) );
ao22f01  g7582 ( .o(n13070), .a(n13069), .b(_net_9242), .c(n10086), .d(_net_9239) );
na02f01  g7583 ( .o(n13071), .a(n13070), .b(n13068) );
ao12f01  g7584 ( .o(n13072), .a(n6490), .b(_net_9244), .c(n8508) );
ao12f01  g7585 ( .o(n13073), .a(n6491), .b(n13072), .c(n6136) );
no04f01  g7586 ( .o(n13074), .a(n13073), .b(n13071), .c(n13067), .d(n13065) );
ao12f01  g7587 ( .o(n6306), .a(n6526_1), .b(n13074), .c(n13064) );
na02f01  g7588 ( .o(n13076), .a(n8841), .b(n10321) );
na02f01  g7589 ( .o(n13077), .a(n5948), .b(net_9251) );
na02f01  g7590 ( .o(n6311), .a(n13077), .b(n13076) );
ao12f01  g7591 ( .o(n13079), .a(n5658), .b(n5678), .c(net_253) );
ao22f01  g7592 ( .o(n13080), .a(n5681_1), .b(x4587), .c(n5680), .d(net_9716) );
na02f01  g7593 ( .o(n6316), .a(n13080), .b(n13079) );
in01f01  g7594 ( .o(n13082), .a(net_10403) );
na02f01  g7595 ( .o(n13083), .a(n8580), .b(net_10385) );
ao12f01  g7596 ( .o(n6321), .a(n11245), .b(n13083), .c(n13082) );
na02f01  g7597 ( .o(n13085), .a(n7937), .b(net_236) );
na02f01  g7598 ( .o(n13086), .a(n7936), .b(net_9766) );
ao22f01  g7599 ( .o(n13087), .a(n7943), .b(_net_10205), .c(n7942), .d(x5790) );
na04f01  g7600 ( .o(n6326), .a(n13087), .b(n13086), .c(n13085), .d(n7939) );
ao12f01  g7601 ( .o(n13089), .a(n5658), .b(n5774), .c(x4781) );
oa12f01  g7602 ( .o(n6331), .a(n13089), .b(n5770), .c(n7027) );
in01f01  g7603 ( .o(n6336), .a(n10152) );
na02f01  g7604 ( .o(n13092), .a(n7353), .b(x5364) );
na02f01  g7605 ( .o(n13093), .a(n7352), .b(net_9674) );
ao22f01  g7606 ( .o(n13094), .a(n7358), .b(net_243), .c(n7357), .d(_net_10107) );
na04f01  g7607 ( .o(n6341), .a(n13094), .b(n13093), .c(n13092), .d(n7355_1) );
na03f01  g7608 ( .o(n13096), .a(n6736), .b(n8525), .c(n12817) );
na04f01  g7609 ( .o(n13097), .a(n6727), .b(n12127), .c(n8661), .d(n6729) );
na04f01  g7610 ( .o(n13098), .a(n10379), .b(n6723_1), .c(n8532), .d(n6720) );
no03f01  g7611 ( .o(n13099), .a(n13098), .b(n13097), .c(n13096) );
ao12f01  g7612 ( .o(n6346), .a(n13099), .b(n11157), .c(n11155) );
in01f01  g7613 ( .o(n13101), .a(net_9504) );
ao22f01  g7614 ( .o(n13102), .a(n5743), .b(x1792), .c(n5742), .d(_net_9413) );
oa12f01  g7615 ( .o(n6351), .a(n13102), .b(n5741), .c(n13101) );
oa22f01  g7616 ( .o(n13104), .a(n6565), .b(n8282), .c(n6563), .d(n12253) );
ao12f01  g7617 ( .o(n13105), .a(n13104), .b(n6555), .c(net_9978) );
ao22f01  g7618 ( .o(n13106), .a(n6573), .b(net_9879), .c(n6572), .d(net_10395) );
ao22f01  g7619 ( .o(n13107), .a(n6580), .b(net_9812), .c(n6577), .d(net_9681) );
na02f01  g7620 ( .o(n13108), .a(n6582), .b(net_9911) );
ao22f01  g7621 ( .o(n13109), .a(n6585), .b(net_9713), .c(n6584_1), .d(net_9780) );
na02f01  g7622 ( .o(n13110), .a(n13109), .b(n13108) );
oa22f01  g7623 ( .o(n13111), .a(n6593), .b(n11803), .c(n6591), .d(n5836) );
oa22f01  g7624 ( .o(n13112), .a(n6600), .b(n5806), .c(n6598), .d(n5778) );
ao22f01  g7625 ( .o(n13113), .a(n6603), .b(net_10500), .c(n6602), .d(net_10010) );
ao22f01  g7626 ( .o(n13114), .a(n6606), .b(_net_9942), .c(n6605), .d(net_10290) );
na02f01  g7627 ( .o(n13115), .a(n13114), .b(n13113) );
no04f01  g7628 ( .o(n13116), .a(n13115), .b(n13112), .c(n13111), .d(n13110) );
na04f01  g7629 ( .o(n6356), .a(n13116), .b(n13107), .c(n13106), .d(n13105) );
no02f01  g7630 ( .o(n6364), .a(n9882), .b(_net_9606) );
in01f01  g7631 ( .o(n13119), .a(net_9946) );
no02f01  g7632 ( .o(n13120), .a(n6973), .b(n9976) );
na03f01  g7633 ( .o(n13121), .a(n5691), .b(x4520), .c(x6599) );
no02f01  g7634 ( .o(n13122), .a(n13120), .b(n5691) );
na02f01  g7635 ( .o(n13123), .a(n13122), .b(x6599) );
oa12f01  g7636 ( .o(n6373), .a(n13121), .b(n13123), .c(n13119) );
oa22f01  g7637 ( .o(n6378), .a(n5694), .b(n6964), .c(n5692), .d(n5600) );
na02f01  g7638 ( .o(n13126), .a(n6936), .b(n6903) );
na02f01  g7639 ( .o(n13127), .a(n6170), .b(_net_10259) );
na03f01  g7640 ( .o(n13128), .a(n13127), .b(n13126), .c(n6175) );
oa12f01  g7641 ( .o(n13129), .a(n6907), .b(n6906), .c(n12801) );
in01f01  g7642 ( .o(n13130), .a(n6907) );
no02f01  g7643 ( .o(n13131), .a(n6906), .b(n12801) );
na02f01  g7644 ( .o(n13132), .a(n13131), .b(n13130) );
na03f01  g7645 ( .o(n13133), .a(n13132), .b(n13129), .c(n6177_1) );
na02f01  g7646 ( .o(n13134), .a(n6168), .b(_net_10259) );
na03f01  g7647 ( .o(n6383), .a(n13134), .b(n13133), .c(n13128) );
in01f01  g7648 ( .o(n13136), .a(n8839_1) );
in01f01  g7649 ( .o(n13137), .a(n8842) );
oa12f01  g7650 ( .o(n13138), .a(n13137), .b(n8843), .c(n13136) );
in01f01  g7651 ( .o(n13139), .a(n8843) );
na03f01  g7652 ( .o(n13140), .a(n13139), .b(n8842), .c(n8839_1) );
na02f01  g7653 ( .o(n6388), .a(n13140), .b(n13138) );
oa22f01  g7654 ( .o(n13142), .a(n6565), .b(n11492), .c(n6563), .d(n8256) );
ao12f01  g7655 ( .o(n13143), .a(n13142), .b(n6584_1), .c(net_9768) );
ao22f01  g7656 ( .o(n13144), .a(n6606), .b(_net_9931), .c(n6602), .d(net_9998) );
ao22f01  g7657 ( .o(n13145), .a(n6597), .b(_net_9733), .c(n6580), .d(net_9800) );
na02f01  g7658 ( .o(n13146), .a(n8042), .b(net_10527) );
na02f01  g7659 ( .o(n13147), .a(n6555), .b(net_9966) );
na02f01  g7660 ( .o(n13148), .a(n6577), .b(net_9669) );
na02f01  g7661 ( .o(n13149), .a(n6585), .b(net_9701) );
na04f01  g7662 ( .o(n13150), .a(n13149), .b(n13148), .c(n13147), .d(n13146) );
ao22f01  g7663 ( .o(n13151), .a(n6599_1), .b(_net_9832), .c(n6590), .d(_net_10030) );
na02f01  g7664 ( .o(n13152), .a(n6573), .b(net_9867) );
na02f01  g7665 ( .o(n13153), .a(n6582), .b(net_9899) );
na03f01  g7666 ( .o(n13154), .a(n13153), .b(n13152), .c(n13151) );
no02f01  g7667 ( .o(n13155), .a(n13154), .b(n13150) );
na04f01  g7668 ( .o(n6393), .a(n13155), .b(n13145), .c(n13144), .d(n13143) );
no02f01  g7669 ( .o(n13157), .a(n6026), .b(n7536) );
ao12f01  g7670 ( .o(n13158), .a(n13157), .b(n6028_1), .c(n5998_1) );
oa12f01  g7671 ( .o(n6397), .a(n13158), .b(n6022), .c(n5989) );
na02f01  g7672 ( .o(n13160), .a(n6056), .b(_net_254) );
na02f01  g7673 ( .o(n13161), .a(n6055), .b(net_9982) );
ao22f01  g7674 ( .o(n13162), .a(n6062_1), .b(x4520), .c(n6060), .d(_net_10433) );
na04f01  g7675 ( .o(n6406), .a(n13162), .b(n13161), .c(n13160), .d(n6058) );
in01f01  g7676 ( .o(n13164), .a(_net_10207) );
ao12f01  g7677 ( .o(n13165), .a(n5658), .b(n6887), .c(x5647) );
oa12f01  g7678 ( .o(n6411), .a(n13165), .b(n6885_1), .c(n13164) );
in01f01  g7679 ( .o(n13167), .a(_net_10427) );
ao12f01  g7680 ( .o(n13168), .a(n5658), .b(n6052_1), .c(x5003) );
oa12f01  g7681 ( .o(n6416), .a(n13168), .b(n6048), .c(n13167) );
na03f01  g7682 ( .o(n13170), .a(_net_10114), .b(_net_10115), .c(_net_10116) );
na02f01  g7683 ( .o(n6421), .a(n13170), .b(n5749) );
no02f01  g7684 ( .o(n13172), .a(n8813), .b(_net_9293) );
na02f01  g7685 ( .o(n13173), .a(n9811), .b(n8809_1) );
oa22f01  g7686 ( .o(n6426), .a(n13173), .b(n13172), .c(n8817), .d(n7073_1) );
ao12f01  g7687 ( .o(n13175), .a(n5658), .b(n6875_1), .c(net_262) );
ao22f01  g7688 ( .o(n13176), .a(n6878), .b(x3889), .c(n6877), .d(net_9923) );
na02f01  g7689 ( .o(n6431), .a(n13176), .b(n13175) );
no03f01  g7690 ( .o(n6436), .a(n12589), .b(n8026_1), .c(n7701) );
in01f01  g7691 ( .o(n13179), .a(_net_10310) );
ao12f01  g7692 ( .o(n13180), .a(n5658), .b(n5774), .c(x5790) );
oa12f01  g7693 ( .o(n6441), .a(n13180), .b(n5770), .c(n13179) );
in01f01  g7694 ( .o(n13182), .a(net_10405) );
na02f01  g7695 ( .o(n13183), .a(_net_9117), .b(net_10385) );
ao12f01  g7696 ( .o(n6446), .a(n11245), .b(n13183), .c(n13182) );
ao22f01  g7697 ( .o(n13185), .a(n5842), .b(net_9708), .c(n5841), .d(net_148) );
na02f01  g7698 ( .o(n13186), .a(n5847), .b(net_10005) );
ao22f01  g7699 ( .o(n13187), .a(n5850), .b(net_9807), .c(n5849_1), .d(net_9906) );
na03f01  g7700 ( .o(n6451), .a(n13187), .b(n13186), .c(n13185) );
ao22f01  g7701 ( .o(n13189), .a(n5702), .b(x2531), .c(n5701), .d(_net_9401) );
oa12f01  g7702 ( .o(n6456), .a(n13189), .b(n5700_1), .c(n10271) );
in01f01  g7703 ( .o(n13191), .a(net_10495) );
oa22f01  g7704 ( .o(n6469), .a(n7467), .b(n5615), .c(n7465_1), .d(n13191) );
ao12f01  g7705 ( .o(n13193), .a(n5658), .b(n7737), .c(net_9349) );
oa12f01  g7706 ( .o(n6474), .a(n13193), .b(n7736), .c(n8643) );
ao12f01  g7707 ( .o(n13195), .a(n5658), .b(n6532), .c(net_240) );
ao22f01  g7708 ( .o(n13196), .a(n6535), .b(x5548), .c(n6534), .d(net_10000) );
na02f01  g7709 ( .o(n6479), .a(n13196), .b(n13195) );
ao12f01  g7710 ( .o(n13198), .a(n5658), .b(n6887), .c(x3949) );
oa12f01  g7711 ( .o(n6484), .a(n13198), .b(n6885_1), .c(n9220) );
in01f01  g7712 ( .o(n13200), .a(_net_10215) );
ao12f01  g7713 ( .o(n13201), .a(n5658), .b(n6887), .c(x5143) );
oa12f01  g7714 ( .o(n6489), .a(n13201), .b(n6885_1), .c(n13200) );
ao12f01  g7715 ( .o(n13203), .a(n5658), .b(n7844), .c(net_241) );
ao22f01  g7716 ( .o(n13204), .a(n7847), .b(x5498), .c(n7846), .d(net_9803) );
na02f01  g7717 ( .o(n6498), .a(n13204), .b(n13203) );
in01f01  g7718 ( .o(n13206), .a(_net_10111) );
ao12f01  g7719 ( .o(n13207), .a(n5658), .b(n6160_1), .c(x5077) );
oa12f01  g7720 ( .o(n6503), .a(n13207), .b(n6159), .c(n13206) );
oa12f01  g7721 ( .o(n13209), .a(n5880), .b(n5878_1), .c(n5858_1) );
na02f01  g7722 ( .o(n13210), .a(n13209), .b(n5875) );
oa12f01  g7723 ( .o(n13211), .a(n9956), .b(net_9531), .c(net_9542) );
ao12f01  g7724 ( .o(n13212), .a(n5886), .b(n13211), .c(n8399_1) );
ao12f01  g7725 ( .o(n13213), .a(_net_9250), .b(net_9531), .c(n8405) );
no02f01  g7726 ( .o(n13214), .a(n13213), .b(n5891) );
no02f01  g7727 ( .o(n13215), .a(net_9531), .b(_net_9437) );
oa12f01  g7728 ( .o(n13216), .a(x6599), .b(n13215), .c(n13050) );
no03f01  g7729 ( .o(n13217), .a(n13216), .b(n13214), .c(n13212) );
no02f01  g7730 ( .o(n13218), .a(n5858_1), .b(n5658) );
oa12f01  g7731 ( .o(n13219), .a(n8399_1), .b(n5858_1), .c(_net_9437) );
ao22f01  g7732 ( .o(n13220), .a(n13219), .b(n8412), .c(n13218), .d(n5857) );
na03f01  g7733 ( .o(n6512), .a(n13220), .b(n13217), .c(n13210) );
ao22f01  g7734 ( .o(n13222), .a(n5702), .b(x2400), .c(n5701), .d(_net_9403) );
oa12f01  g7735 ( .o(n6517), .a(n13222), .b(n5700_1), .c(n8805) );
in01f01  g7736 ( .o(n13224), .a(x637) );
na02f01  g7737 ( .o(n13225), .a(n10171), .b(n7110) );
na02f01  g7738 ( .o(n13226), .a(n10169), .b(n10326) );
in01f01  g7739 ( .o(n13227), .a(n10174) );
ao22f01  g7740 ( .o(n13228), .a(n10179), .b(n10159), .c(n13227), .d(n10172) );
na03f01  g7741 ( .o(n13229), .a(n13228), .b(n13226), .c(n13225) );
ao12f01  g7742 ( .o(n13230), .a(n13229), .b(n10163), .c(n7140) );
oa22f01  g7743 ( .o(n6522), .a(n13230), .b(n10157), .c(n10155), .d(n13224) );
in01f01  g7744 ( .o(n13232), .a(net_9742) );
oa22f01  g7745 ( .o(n6526), .a(n7367), .b(n13232), .c(n7365_1), .d(n5591) );
ao12f01  g7746 ( .o(n13234), .a(n5658), .b(n5774), .c(x4449) );
oa12f01  g7747 ( .o(n6531), .a(n13234), .b(n5770), .c(n7042) );
ao22f01  g7748 ( .o(n13236), .a(n5842), .b(net_9685), .c(n5841), .d(_net_123) );
na02f01  g7749 ( .o(n13237), .a(n5847), .b(net_9982) );
ao22f01  g7750 ( .o(n13238), .a(n5850), .b(net_9784), .c(n5849_1), .d(net_9883) );
na03f01  g7751 ( .o(n6536), .a(n13238), .b(n13237), .c(n13236) );
na03f01  g7752 ( .o(n13240), .a(n6850), .b(n6486), .c(_net_9235) );
na02f01  g7753 ( .o(n13241), .a(n6471), .b(_net_9235) );
no02f01  g7754 ( .o(n13242), .a(n13241), .b(n7862_1) );
ao12f01  g7755 ( .o(n13243), .a(n6526_1), .b(n10086), .c(_net_9235) );
oa12f01  g7756 ( .o(n13244), .a(n13243), .b(n6477), .c(n10424) );
no02f01  g7757 ( .o(n13245), .a(n13241), .b(n7863) );
no03f01  g7758 ( .o(n13246), .a(n6861_1), .b(n10424), .c(n6511) );
no04f01  g7759 ( .o(n13247), .a(n13246), .b(n13245), .c(n13244), .d(n13242) );
no03f01  g7760 ( .o(n13248), .a(n6474_1), .b(n10424), .c(n6463) );
no02f01  g7761 ( .o(n13249), .a(n6499), .b(n10424) );
oa22f01  g7762 ( .o(n13250), .a(n13241), .b(n7852), .c(n6493_1), .d(n10424) );
no03f01  g7763 ( .o(n13251), .a(n13250), .b(n13249), .c(n13248) );
na03f01  g7764 ( .o(n6541), .a(n13251), .b(n13247), .c(n13240) );
ao22f01  g7765 ( .o(n13253), .a(n5842), .b(net_9680), .c(n5841), .d(_net_118) );
na02f01  g7766 ( .o(n13254), .a(n5847), .b(net_9977) );
ao22f01  g7767 ( .o(n13255), .a(n5850), .b(net_9779), .c(n5849_1), .d(net_9878) );
na03f01  g7768 ( .o(n6546), .a(n13255), .b(n13254), .c(n13253) );
na02f01  g7769 ( .o(n13257), .a(n6056), .b(net_241) );
na02f01  g7770 ( .o(n13258), .a(n6055), .b(net_9969) );
ao22f01  g7771 ( .o(n13259), .a(n6062_1), .b(x5498), .c(n6060), .d(_net_10420) );
na04f01  g7772 ( .o(n6551), .a(n13259), .b(n13258), .c(n13257), .d(n6058) );
ao12f01  g7773 ( .o(n13261), .a(n6131_1), .b(n6148), .c(net_9368) );
oa12f01  g7774 ( .o(n6556), .a(n13261), .b(n8101_1), .c(n7089) );
in01f01  g7775 ( .o(n13263), .a(net_10069) );
in01f01  g7776 ( .o(n13264), .a(net_9659) );
na02f01  g7777 ( .o(n13265), .a(n13264), .b(_net_9660) );
ao12f01  g7778 ( .o(n6561), .a(n6155_1), .b(n13265), .c(n13263) );
na02f01  g7779 ( .o(n13267), .a(n6704_1), .b(n7651) );
na02f01  g7780 ( .o(n13268), .a(n13267), .b(n7653) );
oa22f01  g7781 ( .o(n6566), .a(n13268), .b(n6688), .c(n6685), .d(n7651) );
no02f01  g7782 ( .o(n13270), .a(n6561_1), .b(n10364) );
ao22f01  g7783 ( .o(n13271), .a(n13270), .b(n6558), .c(n6577), .d(net_9691) );
ao22f01  g7784 ( .o(n13272), .a(n6606), .b(net_9952), .c(n6582), .d(net_9921) );
ao22f01  g7785 ( .o(n13273), .a(n6603), .b(net_10496), .c(n6572), .d(net_10391) );
na02f01  g7786 ( .o(n13274), .a(n6580), .b(net_9822) );
ao22f01  g7787 ( .o(n13275), .a(n6605), .b(net_10286), .c(n6585), .d(net_9723) );
na02f01  g7788 ( .o(n13276), .a(n13275), .b(n13274) );
na02f01  g7789 ( .o(n13277), .a(n6555), .b(net_9988) );
na02f01  g7790 ( .o(n13278), .a(n6573), .b(net_9889) );
ao22f01  g7791 ( .o(n13279), .a(n6592), .b(net_10181), .c(n6584_1), .d(net_9790) );
na03f01  g7792 ( .o(n13280), .a(n13279), .b(n13278), .c(n13277) );
ao22f01  g7793 ( .o(n13281), .a(n6602), .b(net_10020), .c(n6599_1), .d(net_9853) );
ao22f01  g7794 ( .o(n13282), .a(n6597), .b(net_9754), .c(n6590), .d(net_10051) );
na02f01  g7795 ( .o(n13283), .a(n13282), .b(n13281) );
no03f01  g7796 ( .o(n13284), .a(n13283), .b(n13280), .c(n13276) );
na04f01  g7797 ( .o(n6571), .a(n13284), .b(n13273), .c(n13272), .d(n13271) );
na02f01  g7798 ( .o(n13286), .a(n7937), .b(net_247) );
na02f01  g7799 ( .o(n13287), .a(n7936), .b(net_9777) );
ao22f01  g7800 ( .o(n13288), .a(n7943), .b(_net_10216), .c(n7942), .d(x5077) );
na04f01  g7801 ( .o(n6575), .a(n13288), .b(n13287), .c(n13286), .d(n7939) );
na02f01  g7802 ( .o(n13290), .a(_net_9606), .b(net_116) );
no02f01  g7803 ( .o(n13291), .a(n7637), .b(n7630) );
oa12f01  g7804 ( .o(n13292), .a(n13291), .b(n7624), .c(n7541) );
in01f01  g7805 ( .o(n13293), .a(n7510) );
no03f01  g7806 ( .o(n13294), .a(n13293), .b(n7625), .c(n7630) );
in01f01  g7807 ( .o(n13295), .a(n13294) );
ao12f01  g7808 ( .o(n13296), .a(_net_9561), .b(n13295), .c(n13292) );
in01f01  g7809 ( .o(n13297), .a(_net_9561) );
in01f01  g7810 ( .o(n13298), .a(n13291) );
ao12f01  g7811 ( .o(n13299), .a(n13298), .b(n7636_1), .c(n10564) );
no03f01  g7812 ( .o(n13300), .a(n13294), .b(n13299), .c(n13297) );
oa12f01  g7813 ( .o(n13301), .a(n7500), .b(n13300), .c(n13296) );
na02f01  g7814 ( .o(n6584), .a(n13301), .b(n13290) );
ao12f01  g7815 ( .o(n13303), .a(n5658), .b(n7844), .c(net_250) );
ao22f01  g7816 ( .o(n13304), .a(n7847), .b(x4851), .c(n7846), .d(net_9812) );
na02f01  g7817 ( .o(n6589), .a(n13304), .b(n13303) );
na03f01  g7818 ( .o(n13306), .a(n5916), .b(n5983_1), .c(n7592) );
na04f01  g7819 ( .o(n13307), .a(n8466), .b(n7554), .c(n8468), .d(n5975) );
na04f01  g7820 ( .o(n13308), .a(n7573), .b(n7071), .c(n5990), .d(n5989) );
no04f01  g7821 ( .o(n6594), .a(n13308), .b(n13307), .c(n13306), .d(n7976) );
na02f01  g7822 ( .o(n13310), .a(n6038), .b(net_235) );
na02f01  g7823 ( .o(n13311), .a(n6037_1), .b(net_9864) );
ao22f01  g7824 ( .o(n13312), .a(n6044), .b(x5850), .c(n6042_1), .d(_net_10309) );
na04f01  g7825 ( .o(n6599), .a(n13312), .b(n13311), .c(n13310), .d(n6040) );
na02f01  g7826 ( .o(n13314), .a(n6349), .b(n6238) );
oa22f01  g7827 ( .o(n6604), .a(n13314), .b(n6348), .c(n6349), .d(n8903) );
in01f01  g7828 ( .o(n13316), .a(net_9753) );
oa12f01  g7829 ( .o(n13317), .a(x6599), .b(n8828), .c(n5674) );
na02f01  g7830 ( .o(n13318), .a(n8830), .b(net_10175) );
oa22f01  g7831 ( .o(n6609), .a(n13318), .b(n8827), .c(n13317), .d(n13316) );
no02f01  g7832 ( .o(n13320), .a(n9914), .b(net_9223) );
no03f01  g7833 ( .o(n6614), .a(n13320), .b(n9916), .c(n9904) );
na04f01  g7834 ( .o(n13322), .a(n10366), .b(n10368), .c(net_9271), .d(x6599) );
oa12f01  g7835 ( .o(n6619), .a(n13322), .b(n10373), .c(n10368) );
in01f01  g7836 ( .o(n13324), .a(n7381) );
na02f01  g7837 ( .o(n13325), .a(n13324), .b(n7419) );
no02f01  g7838 ( .o(n13326), .a(n13325), .b(n7409) );
no02f01  g7839 ( .o(n13327), .a(n7383), .b(n7378) );
in01f01  g7840 ( .o(n13328), .a(n13327) );
ao12f01  g7841 ( .o(n13329), .a(n7875), .b(n13328), .c(n13326) );
oa12f01  g7842 ( .o(n13330), .a(n13329), .b(n13328), .c(n13326) );
na02f01  g7843 ( .o(n13331), .a(n7443), .b(_net_10474) );
na02f01  g7844 ( .o(n13332), .a(n13331), .b(n11567) );
ao22f01  g7845 ( .o(n13333), .a(n13332), .b(n7450), .c(n7453), .d(_net_10474) );
na02f01  g7846 ( .o(n6624), .a(n13333), .b(n13330) );
ao22f01  g7847 ( .o(n13335), .a(n5842), .b(_net_9752), .c(n5841), .d(_net_188) );
na02f01  g7848 ( .o(n13336), .a(n5847), .b(_net_10049) );
ao22f01  g7849 ( .o(n13337), .a(n5850), .b(_net_9851), .c(n5849_1), .d(_net_9950) );
na03f01  g7850 ( .o(n6629), .a(n13337), .b(n13336), .c(n13335) );
in01f01  g7851 ( .o(n13339), .a(n8473) );
oa22f01  g7852 ( .o(n13340), .a(n5916), .b(_net_9291), .c(_net_9290), .d(n7592) );
ao12f01  g7853 ( .o(n13341), .a(n8458), .b(n13340), .c(n8460) );
na02f01  g7854 ( .o(n13342), .a(n7573), .b(_net_9292) );
oa12f01  g7855 ( .o(n13343), .a(n10542), .b(n13342), .c(n8456) );
no02f01  g7856 ( .o(n13344), .a(n13343), .b(n13341) );
no03f01  g7857 ( .o(n13345), .a(n13344), .b(n10543), .c(n13339) );
no02f01  g7858 ( .o(n13346), .a(_net_9297), .b(n7554) );
no02f01  g7859 ( .o(n13347), .a(_net_171), .b(n7605_1) );
ao12f01  g7860 ( .o(n13348), .a(n8470), .b(n8476), .c(n13347) );
oa22f01  g7861 ( .o(n13349), .a(n13348), .b(n13339), .c(n13346), .d(n8467_1) );
no02f01  g7862 ( .o(n13350), .a(n13349), .b(n13345) );
no04f01  g7863 ( .o(n13351), .a(n13350), .b(n8489), .c(n8487), .d(n8486_1) );
in01f01  g7864 ( .o(n13352), .a(n8486_1) );
ao12f01  g7865 ( .o(n13353), .a(n8482_1), .b(n13352), .c(n8481) );
no02f01  g7866 ( .o(n13354), .a(n13353), .b(n8489) );
no04f01  g7867 ( .o(n6634), .a(n13354), .b(n13351), .c(n8483), .d(_net_181) );
in01f01  g7868 ( .o(n13356), .a(net_10289) );
oa22f01  g7869 ( .o(n6639), .a(n9353), .b(n5612), .c(n9352), .d(n13356) );
no02f01  g7870 ( .o(n13358), .a(n7764), .b(n7762) );
na02f01  g7871 ( .o(n13359), .a(n13358), .b(n7817) );
in01f01  g7872 ( .o(n13360), .a(n13358) );
oa12f01  g7873 ( .o(n13361), .a(n13360), .b(n7816_1), .c(n7814) );
na02f01  g7874 ( .o(n6644), .a(n13361), .b(n13359) );
oa22f01  g7875 ( .o(n6649), .a(n5907), .b(n7412), .c(n5905), .d(n5618) );
ao22f01  g7876 ( .o(n13364), .a(n5842), .b(net_9719), .c(n5841), .d(_net_159) );
na02f01  g7877 ( .o(n13365), .a(n5847), .b(net_10016) );
ao22f01  g7878 ( .o(n13366), .a(n5850), .b(net_9818), .c(n5849_1), .d(net_9917) );
na03f01  g7879 ( .o(n6654), .a(n13366), .b(n13365), .c(n13364) );
ao12f01  g7880 ( .o(n13368), .a(n5658), .b(n6875_1), .c(net_238) );
ao22f01  g7881 ( .o(n13369), .a(n6878), .b(x5647), .c(n6877), .d(net_9899) );
na02f01  g7882 ( .o(n6659), .a(n13369), .b(n13368) );
in01f01  g7883 ( .o(n13371), .a(n9176) );
ao12f01  g7884 ( .o(n13372), .a(n9179), .b(n9215), .c(n13371) );
no02f01  g7885 ( .o(n13373), .a(_net_10267), .b(n9180) );
no02f01  g7886 ( .o(n13374), .a(n9216), .b(n13373) );
na02f01  g7887 ( .o(n13375), .a(n13374), .b(n13372) );
in01f01  g7888 ( .o(n13376), .a(n13372) );
in01f01  g7889 ( .o(n13377), .a(n13374) );
na02f01  g7890 ( .o(n13378), .a(n13377), .b(n13376) );
na02f01  g7891 ( .o(n6664), .a(n13378), .b(n13375) );
in01f01  g7892 ( .o(n13380), .a(_net_10095) );
ao12f01  g7893 ( .o(n13381), .a(n5658), .b(n6160_1), .c(x6102) );
oa12f01  g7894 ( .o(n6669), .a(n13381), .b(n6159), .c(n13380) );
no02f01  g7895 ( .o(n13383), .a(n7778_1), .b(n6723_1) );
no02f01  g7896 ( .o(n13384), .a(n8132), .b(n13383) );
no02f01  g7897 ( .o(n13385), .a(_net_10155), .b(_net_9731) );
no02f01  g7898 ( .o(n13386), .a(n7769), .b(n6720) );
no02f01  g7899 ( .o(n13387), .a(n13386), .b(n13385) );
in01f01  g7900 ( .o(n13388), .a(n13387) );
ao12f01  g7901 ( .o(n13389), .a(n6746), .b(n13388), .c(n13384) );
oa12f01  g7902 ( .o(n13390), .a(n13389), .b(n13388), .c(n13384) );
oa12f01  g7903 ( .o(n13391), .a(_net_10155), .b(n8141), .c(_net_10154) );
na02f01  g7904 ( .o(n13392), .a(n13391), .b(n8143) );
ao22f01  g7905 ( .o(n13393), .a(n13392), .b(n6750), .c(n6760), .d(_net_10155) );
na02f01  g7906 ( .o(n6674), .a(n13393), .b(n13390) );
na02f01  g7907 ( .o(n13395), .a(n8202), .b(_net_10364) );
na02f01  g7908 ( .o(n13396), .a(n8188), .b(n7024) );
na02f01  g7909 ( .o(n13397), .a(n8187), .b(_net_10364) );
na03f01  g7910 ( .o(n13398), .a(n13397), .b(n13396), .c(n8200_1) );
oa12f01  g7911 ( .o(n13399), .a(n8172), .b(n8167), .c(n8162) );
in01f01  g7912 ( .o(n13400), .a(n8172) );
no02f01  g7913 ( .o(n13401), .a(n8167), .b(n8162) );
na02f01  g7914 ( .o(n13402), .a(n13401), .b(n13400) );
na03f01  g7915 ( .o(n13403), .a(n13402), .b(n13399), .c(n8183) );
na03f01  g7916 ( .o(n6679), .a(n13403), .b(n13398), .c(n13395) );
ao12f01  g7917 ( .o(n13405), .a(n5658), .b(n5678), .c(net_262) );
ao22f01  g7918 ( .o(n13406), .a(n5681_1), .b(x3889), .c(n5680), .d(net_9725) );
na02f01  g7919 ( .o(n6684), .a(n13406), .b(n13405) );
oa22f01  g7920 ( .o(n6689), .a(n8418), .b(n8733), .c(n8417), .d(n5621) );
na02f01  g7921 ( .o(n13409), .a(n8943), .b(_net_10332) );
na02f01  g7922 ( .o(n6694), .a(n13409), .b(n8945) );
oa12f01  g7923 ( .o(n13411), .a(n9363), .b(n9358), .c(_net_10162) );
oa12f01  g7924 ( .o(n13412), .a(n13411), .b(n9359), .c(n9361) );
in01f01  g7925 ( .o(n13413), .a(n13412) );
no02f01  g7926 ( .o(n13414), .a(n9362), .b(n7821_1) );
ao12f01  g7927 ( .o(n13415), .a(n13413), .b(n13414), .c(n7818) );
in01f01  g7928 ( .o(n13416), .a(n13415) );
no02f01  g7929 ( .o(n13417), .a(n6667), .b(n9658) );
no02f01  g7930 ( .o(n13418), .a(_net_10125), .b(_net_10163) );
no02f01  g7931 ( .o(n13419), .a(n13418), .b(n13417) );
na02f01  g7932 ( .o(n13420), .a(n13419), .b(n13416) );
in01f01  g7933 ( .o(n13421), .a(n13419) );
na02f01  g7934 ( .o(n13422), .a(n13421), .b(n13415) );
na02f01  g7935 ( .o(n6699), .a(n13422), .b(n13420) );
ao12f01  g7936 ( .o(n13424), .a(n5658), .b(n7737), .c(net_9348) );
oa12f01  g7937 ( .o(n6704), .a(n13424), .b(n7736), .c(n10342) );
no02f01  g7938 ( .o(n13426), .a(n8877), .b(n8875) );
no02f01  g7939 ( .o(n13427), .a(n5968), .b(n8862_1) );
no02f01  g7940 ( .o(n13428), .a(n8876_1), .b(n13427) );
in01f01  g7941 ( .o(n13429), .a(n13428) );
oa12f01  g7942 ( .o(n13430), .a(n13429), .b(n13426), .c(n8861) );
in01f01  g7943 ( .o(n13431), .a(n13426) );
na03f01  g7944 ( .o(n13432), .a(n13428), .b(n13431), .c(n8863) );
na02f01  g7945 ( .o(n6709), .a(n13432), .b(n13430) );
oa12f01  g7946 ( .o(n13434), .a(_net_152), .b(_net_151), .c(n7592) );
no03f01  g7947 ( .o(n13435), .a(_net_151), .b(n7592), .c(_net_152) );
oa12f01  g7948 ( .o(n13436), .a(n13434), .b(n13435), .c(_net_168) );
ao22f01  g7949 ( .o(n13437), .a(_net_169), .b(n5936), .c(_net_170), .d(n5939_1) );
na03f01  g7950 ( .o(n13438), .a(n7573), .b(_net_153), .c(_net_154) );
na03f01  g7951 ( .o(n13439), .a(n7573), .b(_net_153), .c(n7071) );
na02f01  g7952 ( .o(n13440), .a(n7071), .b(_net_154) );
na03f01  g7953 ( .o(n13441), .a(n13440), .b(n13439), .c(n13438) );
ao12f01  g7954 ( .o(n13442), .a(n13441), .b(n13437), .c(n13436) );
ao22f01  g7955 ( .o(n13443), .a(n5966), .b(_net_172), .c(_net_171), .d(n5963) );
oa22f01  g7956 ( .o(n13444), .a(n8466), .b(_net_157), .c(n7554), .d(_net_158) );
in01f01  g7957 ( .o(n13445), .a(n13444) );
na02f01  g7958 ( .o(n13446), .a(n13445), .b(n13443) );
na03f01  g7959 ( .o(n13447), .a(n8468), .b(n5975), .c(_net_155) );
na03f01  g7960 ( .o(n13448), .a(_net_156), .b(n8468), .c(_net_155) );
ao12f01  g7961 ( .o(n13449), .a(n13444), .b(n13448), .c(n13447) );
no03f01  g7962 ( .o(n13450), .a(n13444), .b(n5966), .c(_net_172) );
na03f01  g7963 ( .o(n13451), .a(n8466), .b(_net_157), .c(_net_158) );
na02f01  g7964 ( .o(n13452), .a(n7554), .b(_net_158) );
na03f01  g7965 ( .o(n13453), .a(n8466), .b(n7554), .c(_net_157) );
na03f01  g7966 ( .o(n13454), .a(n13453), .b(n13452), .c(n13451) );
no03f01  g7967 ( .o(n13455), .a(n13454), .b(n13450), .c(n13449) );
oa12f01  g7968 ( .o(n13456), .a(n13455), .b(n13446), .c(n13442) );
no02f01  g7969 ( .o(n13457), .a(n5983_1), .b(_net_161) );
oa22f01  g7970 ( .o(n13458), .a(_net_159), .b(n5989), .c(n5990), .d(_net_160) );
no02f01  g7971 ( .o(n13459), .a(n13458), .b(n13457) );
no03f01  g7972 ( .o(n13460), .a(n5995), .b(n5991), .c(_net_175) );
no03f01  g7973 ( .o(n13461), .a(n5995), .b(_net_176), .c(_net_175) );
oa22f01  g7974 ( .o(n13462), .a(_net_177), .b(n5984), .c(_net_176), .d(n5991) );
no03f01  g7975 ( .o(n13463), .a(n13462), .b(n13461), .c(n13460) );
no03f01  g7976 ( .o(n13464), .a(_net_164), .b(_net_162), .c(_net_163) );
oa12f01  g7977 ( .o(n13465), .a(n13464), .b(n13463), .c(n13457) );
ao12f01  g7978 ( .o(n6718), .a(n13465), .b(n13459), .c(n13456) );
in01f01  g7979 ( .o(n13467), .a(_net_10243) );
na02f01  g7980 ( .o(n13468), .a(_net_10244), .b(n13467) );
ao12f01  g7981 ( .o(n6723), .a(n5658), .b(n13468), .c(n12650) );
na02f01  g7982 ( .o(n13470), .a(net_10396), .b(net_10404) );
ao22f01  g7983 ( .o(n13471), .a(net_10395), .b(net_10403), .c(net_10405), .d(net_10397) );
ao22f01  g7984 ( .o(n13472), .a(net_10401), .b(net_10394), .c(net_10399), .d(net_10392) );
ao22f01  g7985 ( .o(n13473), .a(net_10395), .b(net_10402), .c(net_10400), .d(net_10393) );
na04f01  g7986 ( .o(n6728), .a(n13473), .b(n13472), .c(n13471), .d(n13470) );
ao22f01  g7987 ( .o(n13475), .a(n5842), .b(net_9706), .c(n5841), .d(net_146) );
na02f01  g7988 ( .o(n13476), .a(n5847), .b(net_10003) );
ao22f01  g7989 ( .o(n13477), .a(n5850), .b(net_9805), .c(n5849_1), .d(net_9904) );
na03f01  g7990 ( .o(n6733), .a(n13477), .b(n13476), .c(n13475) );
oa22f01  g7991 ( .o(n6738), .a(n7467), .b(n5597_1), .c(n7465_1), .d(n8608) );
in01f01  g7992 ( .o(n13480), .a(net_9754) );
oa22f01  g7993 ( .o(n6743), .a(n13318), .b(n10282), .c(n13317), .d(n13480) );
na02f01  g7994 ( .o(n13482), .a(n7913), .b(net_9622) );
ao12f01  g7995 ( .o(n6748), .a(n5658), .b(n13482), .c(n7910) );
na02f01  g7996 ( .o(n13484), .a(n7353), .b(x5790) );
na02f01  g7997 ( .o(n13485), .a(n7352), .b(net_9667) );
ao22f01  g7998 ( .o(n13486), .a(n7358), .b(net_236), .c(n7357), .d(_net_10100) );
na04f01  g7999 ( .o(n6753), .a(n13486), .b(n13485), .c(n13484), .d(n7355_1) );
ao12f01  g8000 ( .o(n13488), .a(n5658), .b(n6160_1), .c(x4285) );
oa12f01  g8001 ( .o(n6758), .a(n13488), .b(n6159), .c(n7807) );
oa12f01  g8002 ( .o(n13490), .a(_net_118), .b(n7592), .c(_net_117) );
no03f01  g8003 ( .o(n13491), .a(_net_118), .b(n7592), .c(_net_117) );
oa12f01  g8004 ( .o(n13492), .a(n13490), .b(n13491), .c(_net_168) );
in01f01  g8005 ( .o(n13493), .a(_net_119) );
in01f01  g8006 ( .o(n13494), .a(_net_120) );
ao22f01  g8007 ( .o(n13495), .a(_net_169), .b(n13493), .c(_net_170), .d(n13494) );
na03f01  g8008 ( .o(n13496), .a(n7573), .b(_net_120), .c(_net_119) );
na03f01  g8009 ( .o(n13497), .a(n7573), .b(n7071), .c(_net_119) );
na02f01  g8010 ( .o(n13498), .a(n7071), .b(_net_120) );
na03f01  g8011 ( .o(n13499), .a(n13498), .b(n13497), .c(n13496) );
ao12f01  g8012 ( .o(n13500), .a(n13499), .b(n13495), .c(n13492) );
in01f01  g8013 ( .o(n13501), .a(_net_122) );
in01f01  g8014 ( .o(n13502), .a(_net_121) );
ao22f01  g8015 ( .o(n13503), .a(_net_171), .b(n13502), .c(_net_172), .d(n13501) );
oa22f01  g8016 ( .o(n13504), .a(n8466), .b(_net_123), .c(n7554), .d(_net_124) );
in01f01  g8017 ( .o(n13505), .a(n13504) );
na02f01  g8018 ( .o(n13506), .a(n13505), .b(n13503) );
na03f01  g8019 ( .o(n13507), .a(n8468), .b(_net_121), .c(n5975) );
na03f01  g8020 ( .o(n13508), .a(n8468), .b(_net_121), .c(_net_122) );
ao12f01  g8021 ( .o(n13509), .a(n13504), .b(n13508), .c(n13507) );
no03f01  g8022 ( .o(n13510), .a(n13504), .b(_net_172), .c(n13501) );
na03f01  g8023 ( .o(n13511), .a(n8466), .b(_net_123), .c(_net_124) );
na02f01  g8024 ( .o(n13512), .a(n7554), .b(_net_124) );
na03f01  g8025 ( .o(n13513), .a(n8466), .b(_net_123), .c(n7554) );
na03f01  g8026 ( .o(n13514), .a(n13513), .b(n13512), .c(n13511) );
no03f01  g8027 ( .o(n13515), .a(n13514), .b(n13510), .c(n13509) );
oa12f01  g8028 ( .o(n13516), .a(n13515), .b(n13506), .c(n13500) );
no02f01  g8029 ( .o(n13517), .a(n5983_1), .b(_net_127) );
oa22f01  g8030 ( .o(n13518), .a(n5990), .b(_net_126), .c(n5989), .d(_net_125) );
no02f01  g8031 ( .o(n13519), .a(n13518), .b(n13517) );
in01f01  g8032 ( .o(n13520), .a(_net_126) );
no02f01  g8033 ( .o(n13521), .a(n13520), .b(_net_175) );
na03f01  g8034 ( .o(n13522), .a(n5990), .b(n5989), .c(_net_125) );
ao22f01  g8035 ( .o(n13523), .a(n5983_1), .b(_net_127), .c(n5990), .d(_net_126) );
na02f01  g8036 ( .o(n13524), .a(n13523), .b(n13522) );
ao12f01  g8037 ( .o(n13525), .a(n13524), .b(n13521), .c(_net_125) );
no03f01  g8038 ( .o(n13526), .a(_net_128), .b(_net_129), .c(_net_130) );
oa12f01  g8039 ( .o(n13527), .a(n13526), .b(n13525), .c(n13517) );
ao12f01  g8040 ( .o(n6763), .a(n13527), .b(n13519), .c(n13516) );
na02f01  g8041 ( .o(n13529), .a(n7937), .b(net_251) );
na02f01  g8042 ( .o(n13530), .a(n7936), .b(net_9781) );
ao22f01  g8043 ( .o(n13531), .a(n7943), .b(_net_10220), .c(n7942), .d(x4781) );
na04f01  g8044 ( .o(n6768), .a(n13531), .b(n13530), .c(n13529), .d(n7939) );
in01f01  g8045 ( .o(n13533), .a(_net_9188) );
oa22f01  g8046 ( .o(n6773), .a(n8349_1), .b(n8021_1), .c(n8347), .d(n13533) );
ao22f01  g8047 ( .o(n13535), .a(n5842), .b(net_9738), .c(n5841), .d(_net_179) );
na02f01  g8048 ( .o(n13536), .a(n5847), .b(net_10035) );
ao22f01  g8049 ( .o(n13537), .a(n5850), .b(net_9837), .c(n5849_1), .d(net_9936) );
na03f01  g8050 ( .o(n6778), .a(n13537), .b(n13536), .c(n13535) );
in01f01  g8051 ( .o(n13539), .a(net_10399) );
na02f01  g8052 ( .o(n13540), .a(n10500), .b(net_10385) );
ao12f01  g8053 ( .o(n6786), .a(n11245), .b(n13540), .c(n13539) );
na02f01  g8054 ( .o(n13542), .a(n7937), .b(_net_261) );
na02f01  g8055 ( .o(n13543), .a(n7936), .b(net_9791) );
ao22f01  g8056 ( .o(n13544), .a(n7943), .b(_net_10230), .c(n7942), .d(x3949) );
na04f01  g8057 ( .o(n6791), .a(n13544), .b(n13543), .c(n13542), .d(n7939) );
na02f01  g8058 ( .o(n13546), .a(n7358), .b(_net_259) );
na02f01  g8059 ( .o(n13547), .a(n7352), .b(net_9690) );
ao22f01  g8060 ( .o(n13548), .a(n7357), .b(_net_10123), .c(n7353), .d(x4117) );
na04f01  g8061 ( .o(n6796), .a(n13548), .b(n13547), .c(n13546), .d(n7355_1) );
na02f01  g8062 ( .o(n13550), .a(n6038), .b(net_236) );
na02f01  g8063 ( .o(n13551), .a(n6037_1), .b(net_9865) );
ao22f01  g8064 ( .o(n13552), .a(n6044), .b(x5790), .c(n6042_1), .d(_net_10310) );
na04f01  g8065 ( .o(n6801), .a(n13552), .b(n13551), .c(n13550), .d(n6040) );
na02f01  g8066 ( .o(n13554), .a(n7937), .b(net_241) );
na02f01  g8067 ( .o(n13555), .a(n7936), .b(net_9771) );
ao22f01  g8068 ( .o(n13556), .a(n7943), .b(_net_10210), .c(n7942), .d(x5498) );
na04f01  g8069 ( .o(n6806), .a(n13556), .b(n13555), .c(n13554), .d(n7939) );
ao22f01  g8070 ( .o(n13558), .a(n5842), .b(_net_9732), .c(n5841), .d(_net_173) );
na02f01  g8071 ( .o(n13559), .a(n5847), .b(_net_10029) );
ao22f01  g8072 ( .o(n13560), .a(n5850), .b(_net_9831), .c(n5849_1), .d(_net_9930) );
na03f01  g8073 ( .o(n6811), .a(n13560), .b(n13559), .c(n13558) );
in01f01  g8074 ( .o(n13562), .a(net_9586) );
no02f01  g8075 ( .o(n6816), .a(n13562), .b(_net_9606) );
oa22f01  g8076 ( .o(n6821), .a(n6989_1), .b(n5640), .c(n6988), .d(n10702) );
oa22f01  g8077 ( .o(n6826), .a(n7480_1), .b(n5797_1), .c(n7478), .d(n5552_1) );
ao12f01  g8078 ( .o(n13566), .a(n5658), .b(n7844), .c(_net_234) );
ao22f01  g8079 ( .o(n13567), .a(n7847), .b(x5901), .c(n7846), .d(net_9796) );
na02f01  g8080 ( .o(n6831), .a(n13567), .b(n13566) );
na02f01  g8081 ( .o(n13569), .a(n6020), .b(n6024) );
oa12f01  g8082 ( .o(n6836), .a(n13569), .b(n6020), .c(n5916) );
ao22f01  g8083 ( .o(n13571), .a(n5842), .b(net_9702), .c(n5841), .d(net_142) );
na02f01  g8084 ( .o(n13572), .a(n5847), .b(net_9999) );
ao22f01  g8085 ( .o(n13573), .a(n5850), .b(net_9801), .c(n5849_1), .d(net_9900) );
na03f01  g8086 ( .o(n6841), .a(n13573), .b(n13572), .c(n13571) );
in01f01  g8087 ( .o(n13575), .a(n7788) );
no02f01  g8088 ( .o(n13576), .a(n7779), .b(n7773_1) );
in01f01  g8089 ( .o(n13577), .a(n13576) );
na02f01  g8090 ( .o(n13578), .a(n13577), .b(n13575) );
na02f01  g8091 ( .o(n13579), .a(n13576), .b(n7788) );
na02f01  g8092 ( .o(n6846), .a(n13579), .b(n13578) );
na02f01  g8093 ( .o(n13581), .a(n7353), .b(x5289) );
na02f01  g8094 ( .o(n13582), .a(n7352), .b(net_9675) );
ao22f01  g8095 ( .o(n13583), .a(n7358), .b(net_244), .c(n7357), .d(_net_10108) );
na04f01  g8096 ( .o(n6851), .a(n13583), .b(n13582), .c(n13581), .d(n7355_1) );
no02f01  g8097 ( .o(n13585), .a(n9816), .b(_net_9297) );
na02f01  g8098 ( .o(n13586), .a(n9819), .b(n8809_1) );
oa22f01  g8099 ( .o(n6856), .a(n13586), .b(n13585), .c(n8817), .d(n7552_1) );
oa22f01  g8100 ( .o(n6861), .a(n7480_1), .b(n11734), .c(n7478), .d(n5637) );
no02f01  g8101 ( .o(n13589), .a(n8529_1), .b(n8134) );
no02f01  g8102 ( .o(n13590), .a(n8523), .b(n8526) );
in01f01  g8103 ( .o(n13591), .a(n13590) );
ao12f01  g8104 ( .o(n13592), .a(n6746), .b(n13591), .c(n13589) );
oa12f01  g8105 ( .o(n13593), .a(n13592), .b(n13591), .c(n13589) );
na02f01  g8106 ( .o(n13594), .a(n8145_1), .b(_net_10157) );
na02f01  g8107 ( .o(n13595), .a(n13594), .b(n8539) );
ao22f01  g8108 ( .o(n13596), .a(n13595), .b(n6750), .c(n6760), .d(_net_10157) );
na02f01  g8109 ( .o(n6870), .a(n13596), .b(n13593) );
na02f01  g8110 ( .o(n13598), .a(n9064), .b(_net_10222) );
na02f01  g8111 ( .o(n6875), .a(n13598), .b(n9066) );
na02f01  g8112 ( .o(n13600), .a(n6168), .b(_net_10246) );
na02f01  g8113 ( .o(n13601), .a(n6787), .b(n6829) );
na03f01  g8114 ( .o(n13602), .a(n13601), .b(n6831_1), .c(n6175) );
in01f01  g8115 ( .o(n13603), .a(n6789) );
no02f01  g8116 ( .o(n13604), .a(n6790), .b(n6788) );
na02f01  g8117 ( .o(n13605), .a(n13604), .b(n13603) );
oa12f01  g8118 ( .o(n13606), .a(n6789), .b(n6790), .c(n6788) );
na03f01  g8119 ( .o(n13607), .a(n13606), .b(n13605), .c(n6177_1) );
na03f01  g8120 ( .o(n6880), .a(n13607), .b(n13602), .c(n13600) );
in01f01  g8121 ( .o(n13609), .a(_net_9588) );
na02f01  g8122 ( .o(n13610), .a(n8841), .b(n13609) );
na02f01  g8123 ( .o(n6885), .a(n13610), .b(n6629_1) );
ao12f01  g8124 ( .o(n13612), .a(n5658), .b(n6532), .c(net_244) );
ao22f01  g8125 ( .o(n13613), .a(n6535), .b(x5289), .c(n6534), .d(net_10004) );
na02f01  g8126 ( .o(n6890), .a(n13613), .b(n13612) );
no03f01  g8127 ( .o(n6895), .a(n7742), .b(_net_9173), .c(n7740) );
ao12f01  g8128 ( .o(n13616), .a(n5658), .b(n6052_1), .c(x4041) );
oa12f01  g8129 ( .o(n6900), .a(n13616), .b(n6048), .c(n9041) );
oa22f01  g8130 ( .o(n6905), .a(n5907), .b(n7382), .c(n5905), .d(n5649) );
na02f01  g8131 ( .o(n13619), .a(n7358), .b(_net_232) );
na02f01  g8132 ( .o(n13620), .a(n7352), .b(net_9663) );
ao22f01  g8133 ( .o(n13621), .a(n7357), .b(_net_10096), .c(n7353), .d(x6028) );
na04f01  g8134 ( .o(n6914), .a(n13621), .b(n13620), .c(n13619), .d(n7355_1) );
oa12f01  g8135 ( .o(n13623), .a(n10894), .b(n6139), .c(_net_9384) );
na03f01  g8136 ( .o(n13624), .a(n10045), .b(n6130), .c(_net_9384) );
ao22f01  g8137 ( .o(n13625), .a(n10047), .b(n6143), .c(_net_9386), .d(x6599) );
na03f01  g8138 ( .o(n6919), .a(n13625), .b(n13624), .c(n13623) );
ao12f01  g8139 ( .o(n13627), .a(n5658), .b(n6160_1), .c(x4520) );
oa12f01  g8140 ( .o(n6924), .a(n13627), .b(n6159), .c(n7803) );
no02f01  g8141 ( .o(n13629), .a(n7004), .b(n7000) );
na02f01  g8142 ( .o(n13630), .a(n13629), .b(n7058_1) );
in01f01  g8143 ( .o(n13631), .a(n13629) );
oa12f01  g8144 ( .o(n13632), .a(n13631), .b(n7057), .c(n7055) );
na02f01  g8145 ( .o(n6929), .a(n13632), .b(n13630) );
in01f01  g8146 ( .o(n13634), .a(net_10401) );
na02f01  g8147 ( .o(n13635), .a(net_10385), .b(net_264) );
ao12f01  g8148 ( .o(n6934), .a(n11245), .b(n13635), .c(n13634) );
in01f01  g8149 ( .o(n13637), .a(n12410) );
no03f01  g8150 ( .o(n13638), .a(n12411), .b(n13637), .c(n8241) );
in01f01  g8151 ( .o(n13639), .a(n13638) );
no02f01  g8152 ( .o(n13640), .a(n12412), .b(n12408) );
in01f01  g8153 ( .o(n13641), .a(n13640) );
na02f01  g8154 ( .o(n13642), .a(n13641), .b(n13639) );
na02f01  g8155 ( .o(n13643), .a(n13640), .b(n13638) );
na02f01  g8156 ( .o(n6939), .a(n13643), .b(n13642) );
na03f01  g8157 ( .o(n13645), .a(n5880), .b(n5879), .c(_net_9532) );
no02f01  g8158 ( .o(n13646), .a(n5854), .b(_net_9532) );
no03f01  g8159 ( .o(n13647), .a(n13646), .b(n10356), .c(n5856) );
na02f01  g8160 ( .o(n13648), .a(_net_9532), .b(n8405) );
oa22f01  g8161 ( .o(n13649), .a(n13648), .b(n8404_1), .c(n5871), .d(n5490) );
no02f01  g8162 ( .o(n13650), .a(n13649), .b(n13647) );
no02f01  g8163 ( .o(n13651), .a(n5864), .b(net_9542) );
ao22f01  g8164 ( .o(n13652), .a(n13651), .b(n8401), .c(n8412), .d(n7916) );
na03f01  g8165 ( .o(n6949), .a(n13652), .b(n13650), .c(n13645) );
oa22f01  g8166 ( .o(n13654), .a(n12726), .b(n13263), .c(n6563), .d(n12262) );
ao12f01  g8167 ( .o(n13655), .a(n13654), .b(n6555), .c(net_9985) );
ao22f01  g8168 ( .o(n13656), .a(n6573), .b(net_9886), .c(n6572), .d(net_10388) );
ao22f01  g8169 ( .o(n13657), .a(n6602), .b(net_10017), .c(n6577), .d(net_9688) );
na02f01  g8170 ( .o(n13658), .a(n6584_1), .b(net_9787) );
ao22f01  g8171 ( .o(n13659), .a(n6599_1), .b(_net_9850), .c(n6582), .d(net_9918) );
na02f01  g8172 ( .o(n13660), .a(n13659), .b(n13658) );
ao22f01  g8173 ( .o(n13661), .a(n6592), .b(net_10178), .c(n6590), .d(_net_10048) );
ao22f01  g8174 ( .o(n13662), .a(n6597), .b(_net_9751), .c(n6585), .d(net_9720) );
ao22f01  g8175 ( .o(n13663), .a(n6603), .b(net_10493), .c(n6580), .d(net_9819) );
ao22f01  g8176 ( .o(n13664), .a(n6606), .b(_net_9949), .c(n6605), .d(net_10283) );
na04f01  g8177 ( .o(n13665), .a(n13664), .b(n13663), .c(n13662), .d(n13661) );
no02f01  g8178 ( .o(n13666), .a(n13665), .b(n13660) );
na04f01  g8179 ( .o(n6954), .a(n13666), .b(n13657), .c(n13656), .d(n13655) );
na02f01  g8180 ( .o(n13668), .a(n9894), .b(_net_10229) );
na02f01  g8181 ( .o(n6971), .a(n13668), .b(n10942) );
in01f01  g8182 ( .o(n13670), .a(_net_10208) );
ao12f01  g8183 ( .o(n13671), .a(n5658), .b(n6887), .c(x5601) );
oa12f01  g8184 ( .o(n6976), .a(n13671), .b(n6885_1), .c(n13670) );
na02f01  g8185 ( .o(n13673), .a(_net_10383), .b(_net_10382) );
no02f01  g8186 ( .o(n13674), .a(n13673), .b(n9944) );
in01f01  g8187 ( .o(n13675), .a(_net_10384) );
no02f01  g8188 ( .o(n13676), .a(n9945), .b(n13675) );
no03f01  g8189 ( .o(n13677), .a(n13676), .b(n13674), .c(n9939) );
in01f01  g8190 ( .o(n13678), .a(_net_10407) );
ao12f01  g8191 ( .o(n13679), .a(n5658), .b(_net_10406), .c(n13678) );
na02f01  g8192 ( .o(n13680), .a(n13679), .b(x987) );
oa22f01  g8193 ( .o(n6981), .a(n13680), .b(n13677), .c(n13679), .d(n5658) );
ao12f01  g8194 ( .o(n13682), .a(n5658), .b(n7844), .c(net_258) );
ao22f01  g8195 ( .o(n13683), .a(n7847), .b(x4209), .c(n7846), .d(net_9820) );
na02f01  g8196 ( .o(n6989), .a(n13683), .b(n13682) );
in01f01  g8197 ( .o(n13685), .a(_net_10092) );
ao12f01  g8198 ( .o(n6998), .a(n6155_1), .b(n10694), .c(n13685) );
na02f01  g8199 ( .o(n13687), .a(n6020), .b(n8841) );
oa12f01  g8200 ( .o(n7003), .a(n13687), .b(n6020), .c(n7592) );
no02f01  g8201 ( .o(n13689), .a(_net_10152), .b(_net_9728) );
no02f01  g8202 ( .o(n13690), .a(n13689), .b(n8128) );
ao22f01  g8203 ( .o(n13691), .a(n13690), .b(n10948), .c(n6760), .d(_net_10152) );
oa12f01  g8204 ( .o(n7012), .a(n13691), .b(n10398), .c(_net_10152) );
ao12f01  g8205 ( .o(n13693), .a(n5658), .b(n5774), .c(x4359) );
oa12f01  g8206 ( .o(n7017), .a(n13693), .b(n5770), .c(n7049) );
in01f01  g8207 ( .o(n13695), .a(net_10288) );
oa22f01  g8208 ( .o(n7026), .a(n9353), .b(n5591), .c(n9352), .d(n13695) );
in01f01  g8209 ( .o(n13697), .a(net_10075) );
oa22f01  g8210 ( .o(n7034), .a(n6989_1), .b(n5540), .c(n6988), .d(n13697) );
in01f01  g8211 ( .o(n13699), .a(net_10287) );
oa22f01  g8212 ( .o(n7039), .a(n9353), .b(n5576), .c(n9352), .d(n13699) );
ao12f01  g8213 ( .o(n13701), .a(n5658), .b(n7844), .c(net_236) );
ao22f01  g8214 ( .o(n13702), .a(n7847), .b(x5790), .c(n7846), .d(net_9798) );
na02f01  g8215 ( .o(n7048), .a(n13702), .b(n13701) );
na02f01  g8216 ( .o(n13704), .a(_net_9297), .b(_net_9606) );
oa12f01  g8217 ( .o(n7053), .a(n13704), .b(_net_9606), .c(n9868) );
no02f01  g8218 ( .o(n13706), .a(net_9651), .b(net_9650) );
no03f01  g8219 ( .o(n7058), .a(n13706), .b(n8703), .c(net_9151) );
na02f01  g8220 ( .o(n13708), .a(n12553), .b(net_9276) );
na02f01  g8221 ( .o(n13709), .a(n12552), .b(n12551) );
ao12f01  g8222 ( .o(n7063), .a(n10005), .b(n13709), .c(n13708) );
no02f01  g8223 ( .o(n13711), .a(n9812), .b(_net_9295) );
na02f01  g8224 ( .o(n13712), .a(n9815), .b(n8809_1) );
oa22f01  g8225 ( .o(n7068), .a(n13712), .b(n13711), .c(n8817), .d(n8469) );
na02f01  g8226 ( .o(n13714), .a(n8030), .b(net_9180) );
na02f01  g8227 ( .o(n13715), .a(n8029), .b(n8028) );
na02f01  g8228 ( .o(n7073), .a(n13715), .b(n13714) );
no02f01  g8229 ( .o(n7082), .a(n10632), .b(n6882) );
oa22f01  g8230 ( .o(n7091), .a(n11830), .b(n8686), .c(n11829), .d(n12507) );
ao22f01  g8231 ( .o(n13719), .a(n11503), .b(x1865), .c(n11502), .d(_net_9412) );
oa12f01  g8232 ( .o(n7104), .a(n13719), .b(n11501), .c(n9409) );
na02f01  g8233 ( .o(n13721), .a(n7937), .b(net_248) );
na02f01  g8234 ( .o(n13722), .a(n7936), .b(net_9778) );
ao22f01  g8235 ( .o(n13723), .a(n7943), .b(_net_10217), .c(n7942), .d(x5003) );
na04f01  g8236 ( .o(n7113), .a(n13723), .b(n13722), .c(n13721), .d(n7939) );
oa22f01  g8237 ( .o(n7118), .a(n5907), .b(n5836), .c(n5905), .d(n5546) );
na02f01  g8238 ( .o(n13726), .a(n7937), .b(_net_259) );
na02f01  g8239 ( .o(n13727), .a(n7936), .b(net_9789) );
ao22f01  g8240 ( .o(n13728), .a(n7943), .b(_net_10228), .c(n7942), .d(x4117) );
na04f01  g8241 ( .o(n7123), .a(n13728), .b(n13727), .c(n13726), .d(n7939) );
ao12f01  g8242 ( .o(n13730), .a(n5658), .b(n6052_1), .c(x4520) );
oa12f01  g8243 ( .o(n7128), .a(n13730), .b(n6048), .c(n8213) );
in01f01  g8244 ( .o(n13732), .a(net_10074) );
oa22f01  g8245 ( .o(n7133), .a(n6989_1), .b(n5621), .c(n6988), .d(n13732) );
in01f01  g8246 ( .o(n13734), .a(_net_10099) );
ao12f01  g8247 ( .o(n13735), .a(n5658), .b(n6160_1), .c(x5850) );
oa12f01  g8248 ( .o(n7138), .a(n13735), .b(n6159), .c(n13734) );
no02f01  g8249 ( .o(n13737), .a(n12407), .b(n12404) );
na02f01  g8250 ( .o(n13738), .a(n13737), .b(n12419) );
in01f01  g8251 ( .o(n13739), .a(n13737) );
oa12f01  g8252 ( .o(n13740), .a(n13739), .b(n12418), .c(n12416) );
na02f01  g8253 ( .o(n7143), .a(n13740), .b(n13738) );
ao12f01  g8254 ( .o(n13742), .a(n5658), .b(n5678), .c(net_241) );
ao22f01  g8255 ( .o(n13743), .a(n5681_1), .b(x5498), .c(n5680), .d(net_9704) );
na02f01  g8256 ( .o(n7148), .a(n13743), .b(n13742) );
ao12f01  g8257 ( .o(n13745), .a(n5658), .b(n7844), .c(net_243) );
ao22f01  g8258 ( .o(n13746), .a(n7847), .b(x5364), .c(n7846), .d(net_9805) );
na02f01  g8259 ( .o(n7153), .a(n13746), .b(n13745) );
no02f01  g8260 ( .o(n13748), .a(n6026), .b(n7516) );
ao12f01  g8261 ( .o(n13749), .a(n13748), .b(n6028_1), .c(n5987) );
oa12f01  g8262 ( .o(n7158), .a(n13749), .b(n6022), .c(n5983_1) );
in01f01  g8263 ( .o(n13751), .a(n8888) );
na02f01  g8264 ( .o(n13752), .a(n13751), .b(n10676) );
na02f01  g8265 ( .o(n13753), .a(n13752), .b(n8905) );
no02f01  g8266 ( .o(n13754), .a(n5993_1), .b(n12482) );
no02f01  g8267 ( .o(n13755), .a(n13754), .b(n8887) );
in01f01  g8268 ( .o(n13756), .a(n13755) );
na02f01  g8269 ( .o(n13757), .a(n13756), .b(n13753) );
na03f01  g8270 ( .o(n13758), .a(n13755), .b(n13752), .c(n8905) );
na02f01  g8271 ( .o(n7163), .a(n13758), .b(n13757) );
no02f01  g8272 ( .o(n13760), .a(n10376), .b(n10375) );
ao12f01  g8273 ( .o(n13761), .a(n6746), .b(n13760), .c(n10388) );
oa12f01  g8274 ( .o(n13762), .a(n13761), .b(n13760), .c(n10388) );
na02f01  g8275 ( .o(n13763), .a(n10394), .b(_net_10160) );
ao12f01  g8276 ( .o(n13764), .a(n10398), .b(n12437), .c(n7763_1) );
ao22f01  g8277 ( .o(n13765), .a(n13764), .b(n13763), .c(n6760), .d(_net_10160) );
na02f01  g8278 ( .o(n7168), .a(n13765), .b(n13762) );
ao22f01  g8279 ( .o(n13767), .a(n8047), .b(net_10065), .c(n6564), .d(net_10087) );
oa12f01  g8280 ( .o(n13768), .a(n13767), .b(n6563), .c(n9577) );
ao22f01  g8281 ( .o(n13769), .a(n6590), .b(net_10044), .c(n6580), .d(net_9815) );
na02f01  g8282 ( .o(n13770), .a(n6584_1), .b(net_9783) );
na02f01  g8283 ( .o(n13771), .a(n6602), .b(net_10013) );
na03f01  g8284 ( .o(n13772), .a(n13771), .b(n13770), .c(n13769) );
no02f01  g8285 ( .o(n13773), .a(n13772), .b(n13768) );
ao22f01  g8286 ( .o(n13774), .a(n6585), .b(net_9716), .c(n6573), .d(net_9882) );
ao22f01  g8287 ( .o(n13775), .a(n6582), .b(net_9914), .c(n6555), .d(net_9981) );
in01f01  g8288 ( .o(n13776), .a(net_9945) );
oa22f01  g8289 ( .o(n13777), .a(n6966_1), .b(n13776), .c(n6598), .d(n11072) );
na02f01  g8290 ( .o(n13778), .a(n6577), .b(net_9684) );
oa12f01  g8291 ( .o(n13779), .a(n13778), .b(n6600), .c(n9825) );
no02f01  g8292 ( .o(n13780), .a(n13779), .b(n13777) );
na04f01  g8293 ( .o(n7173), .a(n13780), .b(n13775), .c(n13774), .d(n13773) );
no02f01  g8294 ( .o(n13782), .a(n9912), .b(net_9222) );
no03f01  g8295 ( .o(n7177), .a(n13782), .b(n9914), .c(n9904) );
in01f01  g8296 ( .o(n13784), .a(net_10389) );
oa22f01  g8297 ( .o(n7182), .a(n10211), .b(n5637), .c(n10210), .d(n13784) );
oa22f01  g8298 ( .o(n7187), .a(n5907), .b(n5827), .c(n5905), .d(n5552_1) );
ao12f01  g8299 ( .o(n13787), .a(n5658), .b(n5678), .c(net_239) );
ao22f01  g8300 ( .o(n13788), .a(n5681_1), .b(x5601), .c(n5680), .d(net_9702) );
na02f01  g8301 ( .o(n7192), .a(n13788), .b(n13787) );
no02f01  g8302 ( .o(n13790), .a(n2794), .b(n7590) );
na02f01  g8303 ( .o(n7197), .a(n13790), .b(n5844_1) );
in01f01  g8304 ( .o(n13792), .a(_net_10200) );
ao12f01  g8305 ( .o(n13793), .a(n5658), .b(n6887), .c(x6102) );
oa12f01  g8306 ( .o(n7202), .a(n13793), .b(n6885_1), .c(n13792) );
na02f01  g8307 ( .o(n13795), .a(n5505), .b(n5494) );
no03f01  g8308 ( .o(n7211), .a(n13795), .b(n5497), .c(n5658) );
in01f01  g8309 ( .o(n13797), .a(net_9855) );
oa22f01  g8310 ( .o(n7216), .a(n12533), .b(n8686), .c(n12532), .d(n13797) );
ao22f01  g8311 ( .o(n13799), .a(n5702), .b(x2767), .c(n5701), .d(_net_9397) );
oa12f01  g8312 ( .o(n7221), .a(n13799), .b(n5700_1), .c(n13101) );
na02f01  g8313 ( .o(n13801), .a(n7923), .b(_net_8824) );
na02f01  g8314 ( .o(n13802), .a(n8756), .b(_net_9352) );
ao12f01  g8315 ( .o(n7226), .a(n5658), .b(n13802), .c(n13801) );
ao22f01  g8316 ( .o(n13804), .a(n6602), .b(net_9997), .c(n6597), .d(_net_9732) );
ao22f01  g8317 ( .o(n13805), .a(n6606), .b(_net_9930), .c(n6573), .d(net_9866) );
in01f01  g8318 ( .o(n13806), .a(net_10078) );
ao22f01  g8319 ( .o(n13807), .a(n8045), .b(net_230), .c(n6562), .d(net_203) );
oa12f01  g8320 ( .o(n13808), .a(n13807), .b(n6565), .c(n13806) );
na02f01  g8321 ( .o(n13809), .a(n6577), .b(net_9668) );
na02f01  g8322 ( .o(n13810), .a(n6584_1), .b(net_9767) );
na02f01  g8323 ( .o(n13811), .a(n13810), .b(n13809) );
no02f01  g8324 ( .o(n13812), .a(n13811), .b(n13808) );
ao22f01  g8325 ( .o(n13813), .a(n6603), .b(net_10510), .c(n6585), .d(net_9700) );
oa12f01  g8326 ( .o(n13814), .a(n13813), .b(n8302), .c(n11633) );
ao22f01  g8327 ( .o(n13815), .a(n6590), .b(_net_10029), .c(n6580), .d(net_9799) );
ao22f01  g8328 ( .o(n13816), .a(n6599_1), .b(_net_9831), .c(n6555), .d(net_9965) );
ao22f01  g8329 ( .o(n13817), .a(n6592), .b(net_10195), .c(n6572), .d(net_10405) );
ao22f01  g8330 ( .o(n13818), .a(n8042), .b(net_10526), .c(n6582), .d(net_9898) );
na04f01  g8331 ( .o(n13819), .a(n13818), .b(n13817), .c(n13816), .d(n13815) );
no02f01  g8332 ( .o(n13820), .a(n13819), .b(n13814) );
na04f01  g8333 ( .o(n7231), .a(n13820), .b(n13812), .c(n13805), .d(n13804) );
in01f01  g8334 ( .o(n13822), .a(net_10035) );
oa22f01  g8335 ( .o(n7235), .a(n5907), .b(n13822), .c(n5905), .d(n5634) );
na02f01  g8336 ( .o(n13824), .a(n7353), .b(x5548) );
na02f01  g8337 ( .o(n13825), .a(n7352), .b(net_9671) );
ao22f01  g8338 ( .o(n13826), .a(n7358), .b(net_240), .c(n7357), .d(_net_10104) );
na04f01  g8339 ( .o(n7240), .a(n13826), .b(n13825), .c(n13824), .d(n7355_1) );
na02f01  g8340 ( .o(n13828), .a(n6038), .b(net_245) );
na02f01  g8341 ( .o(n13829), .a(n6037_1), .b(net_9874) );
ao22f01  g8342 ( .o(n13830), .a(n6044), .b(x5225), .c(n6042_1), .d(_net_10319) );
na04f01  g8343 ( .o(n7245), .a(n13830), .b(n13829), .c(n13828), .d(n6040) );
oa22f01  g8344 ( .o(n7250), .a(n5907), .b(n8621_1), .c(n5905), .d(n5603) );
in01f01  g8345 ( .o(n13833), .a(net_10184) );
oa22f01  g8346 ( .o(n7255), .a(n7956), .b(n5612), .c(n7955), .d(n13833) );
ao22f01  g8347 ( .o(n13835), .a(n5842), .b(net_9758), .c(n5841), .d(_net_8834) );
na02f01  g8348 ( .o(n13836), .a(n5847), .b(_net_10055) );
ao22f01  g8349 ( .o(n13837), .a(n5850), .b(net_9857), .c(n5849_1), .d(net_9956) );
na03f01  g8350 ( .o(n7260), .a(n13837), .b(n13836), .c(n13835) );
na02f01  g8351 ( .o(n13839), .a(n8809_1), .b(n7593) );
oa12f01  g8352 ( .o(n7265), .a(n13839), .b(n8817), .c(n7593) );
na02f01  g8353 ( .o(n13841), .a(n7358), .b(net_262) );
na02f01  g8354 ( .o(n13842), .a(n7352), .b(net_9693) );
ao22f01  g8355 ( .o(n13843), .a(n7357), .b(_net_10126), .c(n7353), .d(x3889) );
na04f01  g8356 ( .o(n7275), .a(n13843), .b(n13842), .c(n13841), .d(n7355_1) );
na02f01  g8357 ( .o(n13845), .a(n7358), .b(net_250) );
na02f01  g8358 ( .o(n13846), .a(n7352), .b(net_9681) );
ao22f01  g8359 ( .o(n13847), .a(n7357), .b(_net_10114), .c(n7353), .d(x4851) );
na04f01  g8360 ( .o(n7280), .a(n13847), .b(n13846), .c(n13845), .d(n7355_1) );
na02f01  g8361 ( .o(n13849), .a(n7937), .b(_net_233) );
na02f01  g8362 ( .o(n13850), .a(n7936), .b(net_9763) );
ao22f01  g8363 ( .o(n13851), .a(n7943), .b(_net_10202), .c(n7942), .d(x5961) );
na04f01  g8364 ( .o(n7285), .a(n13851), .b(n13850), .c(n13849), .d(n7939) );
in01f01  g8365 ( .o(n13853), .a(net_10504) );
na02f01  g8366 ( .o(n13854), .a(n10500), .b(net_10490) );
ao12f01  g8367 ( .o(n7290), .a(n9667), .b(n13854), .c(n13853) );
in01f01  g8368 ( .o(n13856), .a(_net_198) );
no02f01  g8369 ( .o(n13857), .a(_net_198), .b(net_197) );
na02f01  g8370 ( .o(n13858), .a(n8262), .b(n573) );
oa22f01  g8371 ( .o(n7295), .a(n13858), .b(n13857), .c(n8280), .d(n13856) );
no02f01  g8372 ( .o(n13860), .a(n9920), .b(net_9225) );
no03f01  g8373 ( .o(n7300), .a(n13860), .b(n10510), .c(n9904) );
na02f01  g8374 ( .o(n13862), .a(n7003), .b(n7991) );
in01f01  g8375 ( .o(n13863), .a(_net_9516) );
oa12f01  g8376 ( .o(n13864), .a(x6599), .b(n8002), .c(n13863) );
ao12f01  g8377 ( .o(n13865), .a(n13864), .b(n7998), .c(n13863) );
na02f01  g8378 ( .o(n7312), .a(n13865), .b(n13862) );
ao12f01  g8379 ( .o(n13867), .a(n5658), .b(n6052_1), .c(x4209) );
oa12f01  g8380 ( .o(n7321), .a(n13867), .b(n6048), .c(n9044) );
in01f01  g8381 ( .o(n13869), .a(net_10492) );
oa22f01  g8382 ( .o(n7326), .a(n7467), .b(n5567_1), .c(n7465_1), .d(n13869) );
na02f01  g8383 ( .o(n13871), .a(n6056), .b(net_243) );
na02f01  g8384 ( .o(n13872), .a(n6055), .b(net_9971) );
ao22f01  g8385 ( .o(n13873), .a(n6062_1), .b(x5364), .c(n6060), .d(_net_10422) );
na04f01  g8386 ( .o(n7331), .a(n13873), .b(n13872), .c(n13871), .d(n6058) );
in01f01  g8387 ( .o(n13875), .a(net_10282) );
oa22f01  g8388 ( .o(n7336), .a(n9353), .b(n5567_1), .c(n9352), .d(n13875) );
ao22f01  g8389 ( .o(n13877), .a(n5842), .b(_net_9729), .c(n5841), .d(_net_170) );
na02f01  g8390 ( .o(n13878), .a(n5847), .b(_net_10026) );
ao22f01  g8391 ( .o(n13879), .a(n5850), .b(_net_9828), .c(n5849_1), .d(_net_9927) );
na03f01  g8392 ( .o(n7341), .a(n13879), .b(n13878), .c(n13877) );
in01f01  g8393 ( .o(n13881), .a(net_10396) );
oa22f01  g8394 ( .o(n7346), .a(n10211), .b(n5640), .c(n10210), .d(n13881) );
no02f01  g8395 ( .o(n13883), .a(n7802), .b(n7798) );
in01f01  g8396 ( .o(n13884), .a(n13883) );
oa12f01  g8397 ( .o(n13885), .a(n13884), .b(n7804), .c(n7793) );
in01f01  g8398 ( .o(n13886), .a(n7793) );
in01f01  g8399 ( .o(n13887), .a(n7804) );
na03f01  g8400 ( .o(n13888), .a(n13883), .b(n13887), .c(n13886) );
na02f01  g8401 ( .o(n7351), .a(n13888), .b(n13885) );
na02f01  g8402 ( .o(n13890), .a(n6056), .b(net_248) );
na02f01  g8403 ( .o(n13891), .a(n6055), .b(net_9976) );
ao22f01  g8404 ( .o(n13892), .a(n6062_1), .b(x5003), .c(n6060), .d(_net_10427) );
na04f01  g8405 ( .o(n7360), .a(n13892), .b(n13891), .c(n13890), .d(n6058) );
oa22f01  g8406 ( .o(n7370), .a(n8418), .b(n8044), .c(n8417), .d(n5540) );
ao22f01  g8407 ( .o(n13895), .a(n5842), .b(net_9694), .c(n5841), .d(net_134) );
na02f01  g8408 ( .o(n13896), .a(n5847), .b(net_9991) );
ao22f01  g8409 ( .o(n13897), .a(n5850), .b(net_9793), .c(n5849_1), .d(net_9892) );
na03f01  g8410 ( .o(n7375), .a(n13897), .b(n13896), .c(n13895) );
no02f01  g8411 ( .o(n7379), .a(n9904), .b(net_9219) );
no02f01  g8412 ( .o(n7384), .a(n10632), .b(n5670) );
na02f01  g8413 ( .o(n13901), .a(n6056), .b(_net_233) );
na02f01  g8414 ( .o(n13902), .a(n6055), .b(net_9961) );
ao22f01  g8415 ( .o(n13903), .a(n6062_1), .b(x5961), .c(n6060), .d(_net_10412) );
na04f01  g8416 ( .o(n7389), .a(n13903), .b(n13902), .c(n13901), .d(n6058) );
in01f01  g8417 ( .o(n13905), .a(n7601) );
ao12f01  g8418 ( .o(n13906), .a(n13905), .b(n6028_1), .c(n5976) );
oa12f01  g8419 ( .o(n7394), .a(n13906), .b(n6022), .c(n5975) );
na02f01  g8420 ( .o(n13908), .a(n6056), .b(net_257) );
na02f01  g8421 ( .o(n13909), .a(n6055), .b(net_9985) );
ao22f01  g8422 ( .o(n13910), .a(n6062_1), .b(x4285), .c(n6060), .d(_net_10436) );
na04f01  g8423 ( .o(n7403), .a(n13910), .b(n13909), .c(n13908), .d(n6058) );
ao22f01  g8424 ( .o(n13912), .a(n5842), .b(net_9750), .c(n5841), .d(net_186) );
na02f01  g8425 ( .o(n13913), .a(n5847), .b(net_10047) );
ao22f01  g8426 ( .o(n13914), .a(n5850), .b(net_9849), .c(n5849_1), .d(net_9948) );
na03f01  g8427 ( .o(n7408), .a(n13914), .b(n13913), .c(n13912) );
in01f01  g8428 ( .o(n13916), .a(_net_10314) );
ao12f01  g8429 ( .o(n13917), .a(n5658), .b(n5774), .c(x5548) );
oa12f01  g8430 ( .o(n7413), .a(n13917), .b(n5770), .c(n13916) );
na02f01  g8431 ( .o(n13919), .a(n7667), .b(n8213) );
na02f01  g8432 ( .o(n13920), .a(n7668), .b(_net_10433) );
na02f01  g8433 ( .o(n7423), .a(n13920), .b(n13919) );
ao22f01  g8434 ( .o(n13922), .a(n5842), .b(net_9703), .c(n5841), .d(net_143) );
na02f01  g8435 ( .o(n13923), .a(n5847), .b(net_10000) );
ao22f01  g8436 ( .o(n13924), .a(n5850), .b(net_9802), .c(n5849_1), .d(net_9901) );
na03f01  g8437 ( .o(n7428), .a(n13924), .b(n13923), .c(n13922) );
oa12f01  g8438 ( .o(n13926), .a(_net_10477), .b(n12405), .c(n9041) );
oa12f01  g8439 ( .o(n13927), .a(n13926), .b(n12406), .c(_net_10439) );
oa12f01  g8440 ( .o(n13928), .a(n13927), .b(n12423), .c(n12421) );
no02f01  g8441 ( .o(n13929), .a(n8793), .b(n7369) );
no02f01  g8442 ( .o(n13930), .a(_net_10440), .b(_net_10478) );
no02f01  g8443 ( .o(n13931), .a(n13930), .b(n13929) );
na02f01  g8444 ( .o(n13932), .a(n13931), .b(n13928) );
in01f01  g8445 ( .o(n13933), .a(n13928) );
in01f01  g8446 ( .o(n13934), .a(n13931) );
na02f01  g8447 ( .o(n13935), .a(n13934), .b(n13933) );
na02f01  g8448 ( .o(n7432), .a(n13935), .b(n13932) );
no02f01  g8449 ( .o(n13937), .a(n11043), .b(net_9231) );
no03f01  g8450 ( .o(n13938), .a(n7704_1), .b(n11343), .c(n11042) );
no03f01  g8451 ( .o(n7441), .a(n13938), .b(n13937), .c(n7703) );
ao22f01  g8452 ( .o(n13940), .a(n5842), .b(net_9698), .c(n5841), .d(net_138) );
na02f01  g8453 ( .o(n13941), .a(n5847), .b(net_9995) );
ao22f01  g8454 ( .o(n13942), .a(n5850), .b(net_9797), .c(n5849_1), .d(net_9896) );
na03f01  g8455 ( .o(n7451), .a(n13942), .b(n13941), .c(n13940) );
ao12f01  g8456 ( .o(n13944), .a(n5658), .b(n6887), .c(x4117) );
oa12f01  g8457 ( .o(n7455), .a(n13944), .b(n6885_1), .c(n9172) );
na02f01  g8458 ( .o(n13946), .a(n6056), .b(_net_259) );
na02f01  g8459 ( .o(n13947), .a(n6055), .b(net_9987) );
ao22f01  g8460 ( .o(n13948), .a(n6062_1), .b(x4117), .c(n6060), .d(_net_10438) );
na04f01  g8461 ( .o(n7460), .a(n13948), .b(n13947), .c(n13946), .d(n6058) );
na02f01  g8462 ( .o(n13950), .a(n8262), .b(n8261) );
na03f01  g8463 ( .o(n13951), .a(n13950), .b(n8264_1), .c(n573) );
oa12f01  g8464 ( .o(n7465), .a(n13951), .b(n8280), .c(n8261) );
no03f01  g8465 ( .o(n13953), .a(n8880), .b(n8866), .c(n8852) );
no02f01  g8466 ( .o(n13954), .a(n5958), .b(n8853_1) );
no02f01  g8467 ( .o(n13955), .a(n8857_1), .b(n13954) );
na02f01  g8468 ( .o(n13956), .a(n13955), .b(n13953) );
in01f01  g8469 ( .o(n13957), .a(n13953) );
in01f01  g8470 ( .o(n13958), .a(n13955) );
na02f01  g8471 ( .o(n13959), .a(n13958), .b(n13957) );
na02f01  g8472 ( .o(n7470), .a(n13959), .b(n13956) );
na02f01  g8473 ( .o(n13961), .a(n8695), .b(net_9152) );
oa12f01  g8474 ( .o(n7475), .a(n13961), .b(n8695), .c(n6357) );
oa22f01  g8475 ( .o(n7484), .a(n7367), .b(n5792_1), .c(n7365_1), .d(n5552_1) );
na02f01  g8476 ( .o(n13964), .a(n6038), .b(_net_232) );
na02f01  g8477 ( .o(n13965), .a(n6037_1), .b(net_9861) );
ao22f01  g8478 ( .o(n13966), .a(n6044), .b(x6028), .c(n6042_1), .d(_net_10306) );
na04f01  g8479 ( .o(n7494), .a(n13966), .b(n13965), .c(n13964), .d(n6040) );
no02f01  g8480 ( .o(n13968), .a(n9201), .b(n9188) );
in01f01  g8481 ( .o(n13969), .a(n13968) );
na02f01  g8482 ( .o(n13970), .a(n13969), .b(n9190) );
na02f01  g8483 ( .o(n13971), .a(n13968), .b(n9191) );
na02f01  g8484 ( .o(n7499), .a(n13971), .b(n13970) );
in01f01  g8485 ( .o(n13973), .a(net_10076) );
oa22f01  g8486 ( .o(n7504), .a(n6989_1), .b(n5573), .c(n6988), .d(n13973) );
in01f01  g8487 ( .o(n13975), .a(net_10400) );
na02f01  g8488 ( .o(n13976), .a(n8768), .b(net_10385) );
ao12f01  g8489 ( .o(n7509), .a(n11245), .b(n13976), .c(n13975) );
in01f01  g8490 ( .o(n13978), .a(_net_10515) );
in01f01  g8491 ( .o(n13979), .a(net_10071) );
ao12f01  g8492 ( .o(n7514), .a(n6155_1), .b(n13979), .c(n13978) );
ao12f01  g8493 ( .o(n13981), .a(n5658), .b(n6532), .c(net_237) );
ao22f01  g8494 ( .o(n13982), .a(n6535), .b(x5722), .c(n6534), .d(net_9997) );
na02f01  g8495 ( .o(n7519), .a(n13982), .b(n13981) );
in01f01  g8496 ( .o(n13984), .a(net_10500) );
oa22f01  g8497 ( .o(n7524), .a(n7467), .b(n5546), .c(n7465_1), .d(n13984) );
in01f01  g8498 ( .o(n13986), .a(net_10391) );
oa22f01  g8499 ( .o(n7529), .a(n10211), .b(n5525), .c(n10210), .d(n13986) );
no02f01  g8500 ( .o(n13988), .a(n9684), .b(n11520) );
in01f01  g8501 ( .o(n13989), .a(n13988) );
no02f01  g8502 ( .o(n13990), .a(n13989), .b(n9678) );
in01f01  g8503 ( .o(n13991), .a(n13990) );
no02f01  g8504 ( .o(n13992), .a(n13991), .b(n6653) );
no02f01  g8505 ( .o(n13993), .a(n9685), .b(n9670) );
ao12f01  g8506 ( .o(n13994), .a(n13993), .b(n8897), .c(net_9599) );
ao12f01  g8507 ( .o(n13995), .a(n13994), .b(n13988), .c(n9674) );
in01f01  g8508 ( .o(n13996), .a(n13995) );
in01f01  g8509 ( .o(n13997), .a(_net_9600) );
no02f01  g8510 ( .o(n13998), .a(n6017), .b(n13997) );
no02f01  g8511 ( .o(n13999), .a(n8912), .b(_net_9600) );
no02f01  g8512 ( .o(n14000), .a(n13999), .b(n13998) );
in01f01  g8513 ( .o(n14001), .a(n14000) );
oa12f01  g8514 ( .o(n14002), .a(n14001), .b(n13996), .c(n13992) );
no02f01  g8515 ( .o(n14003), .a(n13996), .b(n13992) );
na02f01  g8516 ( .o(n14004), .a(n14000), .b(n14003) );
na02f01  g8517 ( .o(n7534), .a(n14004), .b(n14002) );
no02f01  g8518 ( .o(n14006), .a(n9703), .b(n9701) );
ao12f01  g8519 ( .o(n14007), .a(n7875), .b(n14006), .c(n9715) );
oa12f01  g8520 ( .o(n14008), .a(n14007), .b(n14006), .c(n9715) );
no02f01  g8521 ( .o(n14009), .a(n9730), .b(_net_10459) );
no02f01  g8522 ( .o(n14010), .a(n14009), .b(n12277) );
ao22f01  g8523 ( .o(n14011), .a(n14010), .b(n7450), .c(n7453), .d(_net_10459) );
na02f01  g8524 ( .o(n7543), .a(n14011), .b(n14008) );
in01f01  g8525 ( .o(n14013), .a(x769) );
na02f01  g8526 ( .o(n14014), .a(n10171), .b(n7088) );
in01f01  g8527 ( .o(n14015), .a(net_9367) );
na02f01  g8528 ( .o(n14016), .a(n10169), .b(n14015) );
ao22f01  g8529 ( .o(n14017), .a(n13227), .b(net_9270), .c(n10159), .d(_net_9309) );
na03f01  g8530 ( .o(n14018), .a(n14017), .b(n14016), .c(n14014) );
ao12f01  g8531 ( .o(n14019), .a(n14018), .b(n10163), .c(n7319) );
oa22f01  g8532 ( .o(n7548), .a(n14019), .b(n10157), .c(n10155), .d(n14013) );
na02f01  g8533 ( .o(n14021), .a(n9404), .b(n8089) );
na02f01  g8534 ( .o(n14022), .a(n14021), .b(n11821) );
oa22f01  g8535 ( .o(n7552), .a(n14022), .b(n9397), .c(n9407), .d(n8089) );
na02f01  g8536 ( .o(n14024), .a(_net_10172), .b(_net_10173) );
no02f01  g8537 ( .o(n14025), .a(n14024), .b(n9656) );
in01f01  g8538 ( .o(n14026), .a(_net_10174) );
no02f01  g8539 ( .o(n14027), .a(n9657), .b(n14026) );
no03f01  g8540 ( .o(n14028), .a(n14027), .b(n14025), .c(n6979) );
in01f01  g8541 ( .o(n14029), .a(_net_10197) );
ao12f01  g8542 ( .o(n14030), .a(n5658), .b(n14029), .c(_net_10196) );
na02f01  g8543 ( .o(n14031), .a(n14030), .b(x1029) );
oa22f01  g8544 ( .o(n7562), .a(n14031), .b(n14028), .c(n14030), .d(n5658) );
in01f01  g8545 ( .o(n14033), .a(n11841) );
ao12f01  g8546 ( .o(n14034), .a(n11840), .b(n14033), .c(n11839) );
no02f01  g8547 ( .o(n14035), .a(n14034), .b(n9175) );
na02f01  g8548 ( .o(n14036), .a(n14035), .b(_net_10267) );
in01f01  g8549 ( .o(n14037), .a(n14036) );
oa12f01  g8550 ( .o(n14038), .a(n6177_1), .b(n14035), .c(_net_10267) );
na02f01  g8551 ( .o(n14039), .a(n6945), .b(n9185) );
no02f01  g8552 ( .o(n14040), .a(n14039), .b(_net_10266) );
oa12f01  g8553 ( .o(n14041), .a(n6175), .b(n14040), .c(_net_10267) );
ao12f01  g8554 ( .o(n14042), .a(n14041), .b(n14040), .c(_net_10267) );
ao12f01  g8555 ( .o(n14043), .a(n14042), .b(n6168), .c(_net_10267) );
oa12f01  g8556 ( .o(n7566), .a(n14043), .b(n14038), .c(n14037) );
in01f01  g8557 ( .o(n14045), .a(_net_10306) );
ao12f01  g8558 ( .o(n14046), .a(n5658), .b(n5774), .c(x6028) );
oa12f01  g8559 ( .o(n7571), .a(n14046), .b(n5770), .c(n14045) );
na02f01  g8560 ( .o(n14048), .a(n6038), .b(net_256) );
na02f01  g8561 ( .o(n14049), .a(n6037_1), .b(net_9885) );
ao22f01  g8562 ( .o(n14050), .a(n6044), .b(x4359), .c(n6042_1), .d(_net_10330) );
na04f01  g8563 ( .o(n7585), .a(n14050), .b(n14049), .c(n14048), .d(n6040) );
ao22f01  g8564 ( .o(n14052), .a(n5842), .b(net_9672), .c(n5841), .d(net_110) );
na02f01  g8565 ( .o(n14053), .a(n5847), .b(net_9969) );
ao22f01  g8566 ( .o(n14054), .a(n5850), .b(net_9771), .c(n5849_1), .d(net_9870) );
na03f01  g8567 ( .o(n7595), .a(n14054), .b(n14053), .c(n14052) );
oa22f01  g8568 ( .o(n7600), .a(n7367), .b(n6972), .c(n7365_1), .d(n5603) );
ao22f01  g8569 ( .o(n14057), .a(n5842), .b(net_9667), .c(n5841), .d(net_105) );
na02f01  g8570 ( .o(n14058), .a(n5847), .b(net_9964) );
ao22f01  g8571 ( .o(n14059), .a(n5850), .b(net_9766), .c(n5849_1), .d(net_9865) );
na03f01  g8572 ( .o(n7605), .a(n14059), .b(n14058), .c(n14057) );
ao12f01  g8573 ( .o(n14061), .a(n5658), .b(n5678), .c(net_256) );
ao22f01  g8574 ( .o(n14062), .a(n5681_1), .b(x4359), .c(n5680), .d(net_9719) );
na02f01  g8575 ( .o(n7609), .a(n14062), .b(n14061) );
ao22f01  g8576 ( .o(n14064), .a(n5743), .b(x1503), .c(n5742), .d(_net_9418) );
oa12f01  g8577 ( .o(n7621), .a(n14064), .b(n5741), .c(n8114) );
ao12f01  g8578 ( .o(n14066), .a(n5658), .b(n5774), .c(x4209) );
oa12f01  g8579 ( .o(n7626), .a(n14066), .b(n5770), .c(n6999) );
na02f01  g8580 ( .o(n14068), .a(n10370), .b(n11211) );
na02f01  g8581 ( .o(n14069), .a(n14068), .b(n11213) );
oa22f01  g8582 ( .o(n7631), .a(n14069), .b(n10367), .c(n10373), .d(n11211) );
ao12f01  g8583 ( .o(n14071), .a(n5658), .b(n6875_1), .c(net_249) );
ao22f01  g8584 ( .o(n14072), .a(n6878), .b(x4937), .c(n6877), .d(net_9910) );
na02f01  g8585 ( .o(n7636), .a(n14072), .b(n14071) );
in01f01  g8586 ( .o(n14074), .a(net_10505) );
na02f01  g8587 ( .o(n14075), .a(n8768), .b(net_10490) );
ao12f01  g8588 ( .o(n7645), .a(n9667), .b(n14075), .c(n14074) );
no02f01  g8589 ( .o(n14077), .a(n10870), .b(n7416) );
no02f01  g8590 ( .o(n14078), .a(n7414), .b(n7408_1) );
in01f01  g8591 ( .o(n14079), .a(n14078) );
ao12f01  g8592 ( .o(n14080), .a(n7875), .b(n14079), .c(n14077) );
oa12f01  g8593 ( .o(n14081), .a(n14080), .b(n14079), .c(n14077) );
na02f01  g8594 ( .o(n14082), .a(n7439), .b(_net_10472) );
na02f01  g8595 ( .o(n14083), .a(n14082), .b(n7441_1) );
ao22f01  g8596 ( .o(n14084), .a(n14083), .b(n7450), .c(n7453), .d(_net_10472) );
na02f01  g8597 ( .o(n7650), .a(n14084), .b(n14081) );
oa22f01  g8598 ( .o(n7655), .a(n5694), .b(n5707), .c(n5692), .d(n5621) );
na02f01  g8599 ( .o(n14087), .a(n6697), .b(n6690) );
na02f01  g8600 ( .o(n14088), .a(n14087), .b(n6699_1) );
oa22f01  g8601 ( .o(n7660), .a(n14088), .b(n6688), .c(n6685), .d(n6690) );
oa22f01  g8602 ( .o(n7665), .a(n7480_1), .b(n5803), .c(n7478), .d(n5612) );
no02f01  g8603 ( .o(n14091), .a(n8273), .b(net_205) );
oa12f01  g8604 ( .o(n14092), .a(n573), .b(n8274), .c(n8255_1) );
oa22f01  g8605 ( .o(n7670), .a(n14092), .b(n14091), .c(n8280), .d(n8255_1) );
in01f01  g8606 ( .o(n14094), .a(net_10532) );
oa22f01  g8607 ( .o(n7675), .a(n10629), .b(n14094), .c(n8080), .d(n8077) );
ao12f01  g8608 ( .o(n14096), .a(n5658), .b(n5678), .c(net_246) );
ao22f01  g8609 ( .o(n14097), .a(n5681_1), .b(x5143), .c(n5680), .d(net_9709) );
na02f01  g8610 ( .o(n7680), .a(n14097), .b(n14096) );
oa22f01  g8611 ( .o(n7685), .a(n8690), .b(n11828), .c(n8688_1), .d(n11476) );
ao22f01  g8612 ( .o(n14100), .a(n5842), .b(_net_9736), .c(n5841), .d(_net_177) );
na02f01  g8613 ( .o(n14101), .a(n5847), .b(_net_10033) );
ao22f01  g8614 ( .o(n14102), .a(n5850), .b(_net_9835), .c(n5849_1), .d(_net_9934) );
na03f01  g8615 ( .o(n7690), .a(n14102), .b(n14101), .c(n14100) );
ao12f01  g8616 ( .o(n14104), .a(n6933), .b(n14036), .c(n9221) );
oa12f01  g8617 ( .o(n14105), .a(n14104), .b(n14036), .c(n9221) );
na03f01  g8618 ( .o(n14106), .a(n14040), .b(_net_10268), .c(n9171) );
ao12f01  g8619 ( .o(n14107), .a(_net_10268), .b(n14040), .c(n9171) );
no02f01  g8620 ( .o(n14108), .a(n14107), .b(n6846_1) );
ao22f01  g8621 ( .o(n14109), .a(n14108), .b(n14106), .c(n6168), .d(_net_10268) );
na02f01  g8622 ( .o(n7700), .a(n14109), .b(n14105) );
in01f01  g8623 ( .o(n14111), .a(_net_8826) );
na02f01  g8624 ( .o(n7709), .a(n9764), .b(n14111) );
na02f01  g8625 ( .o(n14113), .a(n9771), .b(net_9151) );
no02f01  g8626 ( .o(n14114), .a(n14113), .b(n9758) );
oa12f01  g8627 ( .o(n14115), .a(n9761), .b(n9756), .c(_net_9353) );
oa12f01  g8628 ( .o(n14116), .a(n9771), .b(n8754), .c(net_9151) );
oa12f01  g8629 ( .o(n14117), .a(n9768), .b(n14116), .c(n7886) );
oa12f01  g8630 ( .o(n14118), .a(x6599), .b(n7734_1), .c(n9771) );
ao12f01  g8631 ( .o(n14119), .a(n14118), .b(n9774), .c(_net_9353) );
na02f01  g8632 ( .o(n14120), .a(n14119), .b(n14117) );
ao12f01  g8633 ( .o(n14121), .a(n14120), .b(n14113), .c(n9766) );
oa12f01  g8634 ( .o(n7714), .a(n14121), .b(n14115), .c(n14114) );
ao22f01  g8635 ( .o(n14123), .a(n8118), .b(x3249), .c(n8117), .d(_net_9389) );
oa12f01  g8636 ( .o(n7719), .a(n14123), .b(n8116_1), .c(n13101) );
na02f01  g8637 ( .o(n14125), .a(n9070), .b(_net_10226) );
na02f01  g8638 ( .o(n7724), .a(n14125), .b(n9072) );
in01f01  g8639 ( .o(n14127), .a(_net_10106) );
ao12f01  g8640 ( .o(n14128), .a(n5658), .b(n6160_1), .c(x5427) );
oa12f01  g8641 ( .o(n7729), .a(n14128), .b(n6159), .c(n14127) );
no03f01  g8642 ( .o(n14130), .a(n10314), .b(n9054), .c(_net_10465) );
oa12f01  g8643 ( .o(n14131), .a(n7431), .b(n10315), .c(_net_10466) );
na03f01  g8644 ( .o(n14132), .a(n11337), .b(_net_10466), .c(_net_10465) );
ao12f01  g8645 ( .o(n14133), .a(n7451_1), .b(n12164), .c(n9054) );
ao22f01  g8646 ( .o(n14134), .a(n14133), .b(n14132), .c(n7453), .d(_net_10466) );
oa12f01  g8647 ( .o(n7738), .a(n14134), .b(n14131), .c(n14130) );
oa22f01  g8648 ( .o(n7743), .a(n7367), .b(n8525), .c(n7365_1), .d(n5618) );
na02f01  g8649 ( .o(n14137), .a(n7674), .b(_net_10437) );
na02f01  g8650 ( .o(n7748), .a(n14137), .b(n7676) );
ao12f01  g8651 ( .o(n14139), .a(n6495), .b(n10613), .c(_net_9172) );
na02f01  g8652 ( .o(n14140), .a(_net_9240), .b(_net_9236) );
oa22f01  g8653 ( .o(n14141), .a(n14140), .b(n6861_1), .c(n6493_1), .d(n6495) );
no02f01  g8654 ( .o(n14142), .a(n14141), .b(n14139) );
na02f01  g8655 ( .o(n14143), .a(n6471), .b(_net_9240) );
oa12f01  g8656 ( .o(n14144), .a(_net_9240), .b(n10086), .c(n6476) );
oa12f01  g8657 ( .o(n14145), .a(n14144), .b(n14143), .c(n7863) );
ao12f01  g8658 ( .o(n14146), .a(n14143), .b(n7862_1), .c(n7852) );
na02f01  g8659 ( .o(n14147), .a(n6486), .b(_net_9240) );
ao12f01  g8660 ( .o(n14148), .a(n6463), .b(n6464_1), .c(n6495) );
na02f01  g8661 ( .o(n14149), .a(n14148), .b(n6473) );
oa12f01  g8662 ( .o(n14150), .a(n14149), .b(n14147), .c(n7482) );
no03f01  g8663 ( .o(n14151), .a(n14150), .b(n14146), .c(n14145) );
ao12f01  g8664 ( .o(n7753), .a(n6526_1), .b(n14151), .c(n14142) );
in01f01  g8665 ( .o(n14153), .a(_net_10453) );
na02f01  g8666 ( .o(n14154), .a(_net_10454), .b(n14153) );
ao12f01  g8667 ( .o(n7758), .a(n5658), .b(n14154), .c(n11793) );
no02f01  g8668 ( .o(n7763), .a(n6164_1), .b(n6741) );
in01f01  g8669 ( .o(n14157), .a(_net_10422) );
ao12f01  g8670 ( .o(n14158), .a(n5658), .b(n6052_1), .c(x5364) );
oa12f01  g8671 ( .o(n7768), .a(n14158), .b(n6048), .c(n14157) );
na02f01  g8672 ( .o(n14160), .a(n7450), .b(n9014) );
no02f01  g8673 ( .o(n14161), .a(n9014), .b(_net_10025) );
oa12f01  g8674 ( .o(n14162), .a(n7431), .b(n14161), .c(n9709) );
na02f01  g8675 ( .o(n14163), .a(n7453), .b(_net_10455) );
na03f01  g8676 ( .o(n7773), .a(n14163), .b(n14162), .c(n14160) );
no02f01  g8677 ( .o(n14165), .a(n10256), .b(n7286) );
no02f01  g8678 ( .o(n14166), .a(n10252), .b(n7263) );
no02f01  g8679 ( .o(n14167), .a(n14166), .b(n14165) );
no02f01  g8680 ( .o(n14168), .a(n14167), .b(n7315) );
na02f01  g8681 ( .o(n14169), .a(n14167), .b(n7315) );
na02f01  g8682 ( .o(n14170), .a(n14169), .b(n6148) );
ao12f01  g8683 ( .o(n14171), .a(n6131_1), .b(n6147), .c(net_9368) );
oa12f01  g8684 ( .o(n7778), .a(n14171), .b(n14170), .c(n14168) );
ao12f01  g8685 ( .o(n14173), .a(n5658), .b(n5774), .c(x4587) );
oa12f01  g8686 ( .o(n7787), .a(n14173), .b(n5770), .c(n7017_1) );
ao22f01  g8687 ( .o(n14175), .a(n6590), .b(net_10024), .c(n6580), .d(net_9794) );
ao22f01  g8688 ( .o(n14176), .a(n6584_1), .b(net_9762), .c(n6582), .d(net_9893) );
ao22f01  g8689 ( .o(n14177), .a(n8047), .b(net_10060), .c(n8045), .d(net_225) );
oa12f01  g8690 ( .o(n14178), .a(n14177), .b(n11108), .c(n6514) );
na02f01  g8691 ( .o(n14179), .a(n8042), .b(net_10521) );
ao22f01  g8692 ( .o(n14180), .a(n6564), .b(net_10073), .c(n6562), .d(_net_198) );
na02f01  g8693 ( .o(n14181), .a(n14180), .b(n14179) );
no02f01  g8694 ( .o(n14182), .a(n14181), .b(n14178) );
ao22f01  g8695 ( .o(n14183), .a(n6585), .b(net_9695), .c(n6573), .d(net_9861) );
ao22f01  g8696 ( .o(n14184), .a(n6605), .b(net_10295), .c(n6592), .d(net_10190) );
na02f01  g8697 ( .o(n14185), .a(n14184), .b(n14183) );
ao22f01  g8698 ( .o(n14186), .a(n6602), .b(net_9992), .c(n6572), .d(net_10400) );
ao22f01  g8699 ( .o(n14187), .a(n6603), .b(net_10505), .c(n6577), .d(net_9663) );
ao22f01  g8700 ( .o(n14188), .a(n6606), .b(net_9925), .c(n6597), .d(net_9727) );
ao22f01  g8701 ( .o(n14189), .a(n6599_1), .b(net_9826), .c(n6555), .d(net_9960) );
na04f01  g8702 ( .o(n14190), .a(n14189), .b(n14188), .c(n14187), .d(n14186) );
no02f01  g8703 ( .o(n14191), .a(n14190), .b(n14185) );
na04f01  g8704 ( .o(n7792), .a(n14191), .b(n14182), .c(n14176), .d(n14175) );
ao12f01  g8705 ( .o(n14193), .a(n6131_1), .b(n6148), .c(net_9365) );
oa12f01  g8706 ( .o(n7796), .a(n14193), .b(n8101_1), .c(n7106) );
in01f01  g8707 ( .o(n14195), .a(net_10298) );
na02f01  g8708 ( .o(n14196), .a(n8580), .b(net_10280) );
ao12f01  g8709 ( .o(n7801), .a(n5911), .b(n14196), .c(n14195) );
no02f01  g8710 ( .o(n14198), .a(n8263), .b(_net_200) );
na02f01  g8711 ( .o(n14199), .a(n8266), .b(n573) );
oa22f01  g8712 ( .o(n7806), .a(n14199), .b(n14198), .c(n8280), .d(n8260_1) );
no02f01  g8713 ( .o(n14201), .a(n6822), .b(n6770) );
oa12f01  g8714 ( .o(n14202), .a(n6177_1), .b(n14201), .c(n11508) );
na02f01  g8715 ( .o(n14203), .a(n6841_1), .b(n6770) );
no02f01  g8716 ( .o(n14204), .a(n6842), .b(n6846_1) );
ao22f01  g8717 ( .o(n14205), .a(n14204), .b(n14203), .c(n6168), .d(_net_10254) );
na02f01  g8718 ( .o(n7811), .a(n14205), .b(n14202) );
oa22f01  g8719 ( .o(n7816), .a(n7367), .b(n6723_1), .c(n7365_1), .d(n5573) );
in01f01  g8720 ( .o(n14208), .a(_net_10423) );
ao12f01  g8721 ( .o(n14209), .a(n5658), .b(n6052_1), .c(x5289) );
oa12f01  g8722 ( .o(n7821), .a(n14209), .b(n6048), .c(n14208) );
na02f01  g8723 ( .o(n14211), .a(n6056), .b(net_246) );
na02f01  g8724 ( .o(n14212), .a(n6055), .b(net_9974) );
ao22f01  g8725 ( .o(n14213), .a(n6062_1), .b(x5143), .c(n6060), .d(_net_10425) );
na04f01  g8726 ( .o(n7826), .a(n14213), .b(n14212), .c(n14211), .d(n6058) );
in01f01  g8727 ( .o(n14215), .a(_net_10415) );
ao12f01  g8728 ( .o(n14216), .a(n5658), .b(n6052_1), .c(x5790) );
oa12f01  g8729 ( .o(n7834), .a(n14216), .b(n6048), .c(n14215) );
ao22f01  g8730 ( .o(n14218), .a(n6602), .b(net_9995), .c(n6590), .d(_net_10027) );
ao22f01  g8731 ( .o(n14219), .a(n6584_1), .b(net_9765), .c(n6580), .d(net_9797) );
in01f01  g8732 ( .o(n14220), .a(net_91) );
oa22f01  g8733 ( .o(n14221), .a(n11108), .b(n14220), .c(n6565), .d(n13973) );
oa22f01  g8734 ( .o(n14222), .a(n8046_1), .b(n8416), .c(n6563), .d(n8259) );
oa22f01  g8735 ( .o(n14223), .a(n6966_1), .b(n5711), .c(n6593), .d(n8575) );
no03f01  g8736 ( .o(n14224), .a(n14223), .b(n14222), .c(n14221) );
ao22f01  g8737 ( .o(n14225), .a(n6597), .b(_net_9730), .c(n6585), .d(net_9698) );
oa12f01  g8738 ( .o(n14226), .a(n14225), .b(n8299), .c(n9665) );
ao22f01  g8739 ( .o(n14227), .a(n6582), .b(net_9896), .c(n6577), .d(net_9666) );
ao22f01  g8740 ( .o(n14228), .a(n8042), .b(net_10524), .c(n6605), .d(net_10298) );
ao22f01  g8741 ( .o(n14229), .a(n6573), .b(net_9864), .c(n6572), .d(net_10403) );
ao22f01  g8742 ( .o(n14230), .a(n6599_1), .b(_net_9829), .c(n6555), .d(net_9963) );
na04f01  g8743 ( .o(n14231), .a(n14230), .b(n14229), .c(n14228), .d(n14227) );
no02f01  g8744 ( .o(n14232), .a(n14231), .b(n14226) );
na04f01  g8745 ( .o(n7839), .a(n14232), .b(n14224), .c(n14219), .d(n14218) );
ao12f01  g8746 ( .o(n14234), .a(n5658), .b(n5678), .c(net_243) );
ao22f01  g8747 ( .o(n14235), .a(n5681_1), .b(x5364), .c(n5680), .d(net_9706) );
na02f01  g8748 ( .o(n7843), .a(n14235), .b(n14234) );
oa22f01  g8749 ( .o(n7848), .a(n10323), .b(n8835), .c(n10322), .d(n6097) );
oa22f01  g8750 ( .o(n14238), .a(n12726), .b(n13979), .c(n6563), .d(n10368) );
ao12f01  g8751 ( .o(n14239), .a(n14238), .b(n6555), .c(net_9987) );
ao22f01  g8752 ( .o(n14240), .a(n6573), .b(net_9888), .c(n6572), .d(net_10390) );
ao22f01  g8753 ( .o(n14241), .a(n6602), .b(net_10019), .c(n6577), .d(net_9690) );
na02f01  g8754 ( .o(n14242), .a(n6582), .b(net_9920) );
ao22f01  g8755 ( .o(n14243), .a(n6585), .b(net_9722), .c(n6584_1), .d(net_9789) );
na02f01  g8756 ( .o(n14244), .a(n14243), .b(n14242) );
oa22f01  g8757 ( .o(n14245), .a(n6593), .b(n8440), .c(n6591), .d(n9531) );
oa22f01  g8758 ( .o(n14246), .a(n6600), .b(n11256), .c(n6598), .d(n13316) );
ao22f01  g8759 ( .o(n14247), .a(n6603), .b(net_10495), .c(n6580), .d(net_9821) );
ao22f01  g8760 ( .o(n14248), .a(n6606), .b(net_9951), .c(n6605), .d(net_10285) );
na02f01  g8761 ( .o(n14249), .a(n14248), .b(n14247) );
no04f01  g8762 ( .o(n14250), .a(n14249), .b(n14246), .c(n14245), .d(n14244) );
na04f01  g8763 ( .o(n7853), .a(n14250), .b(n14241), .c(n14240), .d(n14239) );
ao12f01  g8764 ( .o(n14252), .a(n7883), .b(n7923), .c(_net_9313) );
oa12f01  g8765 ( .o(n7857), .a(n14252), .b(n7925_1), .c(n8763) );
na02f01  g8766 ( .o(n14254), .a(n11417), .b(n7902_1) );
na04f01  g8767 ( .o(n14255), .a(n11451), .b(n11421), .c(n5918), .d(_net_185) );
oa12f01  g8768 ( .o(n14256), .a(n11423), .b(n11460), .c(net_9622) );
na03f01  g8769 ( .o(n7866), .a(n14256), .b(n14255), .c(n14254) );
oa22f01  g8770 ( .o(n7871), .a(n7367), .b(n6736), .c(n7365_1), .d(n5561) );
na02f01  g8771 ( .o(n14259), .a(n7423_1), .b(n7371) );
na03f01  g8772 ( .o(n14260), .a(n14259), .b(n7431), .c(n7425) );
no02f01  g8773 ( .o(n14261), .a(n7445), .b(n7371) );
ao12f01  g8774 ( .o(n14262), .a(_net_10476), .b(n7444), .c(n7373) );
no03f01  g8775 ( .o(n14263), .a(n14262), .b(n14261), .c(n7451_1) );
ao12f01  g8776 ( .o(n14264), .a(n14263), .b(n7453), .c(_net_10476) );
na02f01  g8777 ( .o(n7876), .a(n14264), .b(n14260) );
ao12f01  g8778 ( .o(n14266), .a(n5658), .b(n7844), .c(_net_255) );
ao22f01  g8779 ( .o(n14267), .a(n7847), .b(x4449), .c(n7846), .d(net_9817) );
na02f01  g8780 ( .o(n7881), .a(n14267), .b(n14266) );
ao22f01  g8781 ( .o(n14269), .a(n5842), .b(net_9677), .c(n5841), .d(net_115) );
na02f01  g8782 ( .o(n14270), .a(n5847), .b(net_9974) );
ao22f01  g8783 ( .o(n14271), .a(n5850), .b(net_9776), .c(n5849_1), .d(net_9875) );
na03f01  g8784 ( .o(n7889), .a(n14271), .b(n14270), .c(n14269) );
in01f01  g8785 ( .o(n14273), .a(n7615) );
no02f01  g8786 ( .o(n14274), .a(n14273), .b(n7609_1) );
na03f01  g8787 ( .o(n14275), .a(n14274), .b(n7597), .c(n7580_1) );
in01f01  g8788 ( .o(n14276), .a(n14274) );
oa12f01  g8789 ( .o(n14277), .a(n14276), .b(n7633), .c(n7579) );
na02f01  g8790 ( .o(n7893), .a(n14277), .b(n14275) );
in01f01  g8791 ( .o(n14279), .a(net_9925) );
oa22f01  g8792 ( .o(n7898), .a(n5694), .b(n14279), .c(n5692), .d(n5513_1) );
na02f01  g8793 ( .o(n14281), .a(n6038), .b(net_246) );
na02f01  g8794 ( .o(n14282), .a(n6037_1), .b(net_9875) );
ao22f01  g8795 ( .o(n14283), .a(n6044), .b(x5143), .c(n6042_1), .d(_net_10320) );
na04f01  g8796 ( .o(n7911), .a(n14283), .b(n14282), .c(n14281), .d(n6040) );
oa22f01  g8797 ( .o(n14285), .a(n7396), .b(_net_10479), .c(_net_8840), .d(n7399) );
na02f01  g8798 ( .o(n14286), .a(n7396), .b(_net_10479) );
oa22f01  g8799 ( .o(n14287), .a(n7871_1), .b(_net_10481), .c(n7389_1), .d(_net_10480) );
ao12f01  g8800 ( .o(n14288), .a(n14287), .b(n14286), .c(n14285) );
in01f01  g8801 ( .o(n14289), .a(_net_10481) );
oa12f01  g8802 ( .o(n14290), .a(_net_10480), .b(n7871_1), .c(_net_10481) );
oa22f01  g8803 ( .o(n14291), .a(n14290), .b(_net_10027), .c(_net_10028), .d(n14289) );
no02f01  g8804 ( .o(n14292), .a(n14291), .b(n14288) );
oa22f01  g8805 ( .o(n14293), .a(net_10485), .b(n7382), .c(n7379_1), .d(net_10484) );
oa22f01  g8806 ( .o(n14294), .a(n7412), .b(_net_10483), .c(_net_10482), .d(n5897) );
no03f01  g8807 ( .o(n14295), .a(n14294), .b(n14293), .c(n14292) );
in01f01  g8808 ( .o(n14296), .a(_net_10483) );
in01f01  g8809 ( .o(n14297), .a(_net_10482) );
ao12f01  g8810 ( .o(n14298), .a(n14297), .b(_net_10030), .c(n14296) );
ao22f01  g8811 ( .o(n14299), .a(n14298), .b(n5897), .c(n7412), .d(_net_10483) );
oa12f01  g8812 ( .o(n14300), .a(net_10484), .b(net_10485), .c(n7382) );
no02f01  g8813 ( .o(n14301), .a(n14300), .b(_net_10031) );
ao12f01  g8814 ( .o(n14302), .a(n14301), .b(net_10485), .c(n7382) );
oa12f01  g8815 ( .o(n14303), .a(n14302), .b(n14299), .c(n14293) );
oa22f01  g8816 ( .o(n14304), .a(n14303), .b(n14295), .c(_net_10486), .d(n7372) );
na02f01  g8817 ( .o(n14305), .a(_net_10486), .b(n7372) );
no03f01  g8818 ( .o(n14306), .a(net_8835), .b(_net_8821), .c(net_8820) );
na03f01  g8819 ( .o(n7921), .a(n14306), .b(n14305), .c(n14304) );
oa22f01  g8820 ( .o(n7930), .a(n5907), .b(n10292), .c(n5905), .d(n5513_1) );
ao12f01  g8821 ( .o(n14309), .a(n5658), .b(n6532), .c(net_252) );
ao22f01  g8822 ( .o(n14310), .a(n6535), .b(x4694), .c(n6534), .d(net_10012) );
na02f01  g8823 ( .o(n7935), .a(n14310), .b(n14309) );
oa22f01  g8824 ( .o(n7940), .a(n6989_1), .b(n5561), .c(n6988), .d(n13806) );
no02f01  g8825 ( .o(n7945), .a(n7887), .b(n9767) );
oa22f01  g8826 ( .o(n14314), .a(n6600), .b(n6773_1), .c(n6563), .d(n9448) );
na02f01  g8827 ( .o(n14315), .a(n6584_1), .b(net_9771) );
na02f01  g8828 ( .o(n14316), .a(n6573), .b(net_9870) );
ao22f01  g8829 ( .o(n14317), .a(n6597), .b(_net_9736), .c(n6555), .d(net_9969) );
na03f01  g8830 ( .o(n14318), .a(n14317), .b(n14316), .c(n14315) );
no02f01  g8831 ( .o(n14319), .a(n14318), .b(n14314) );
in01f01  g8832 ( .o(n14320), .a(net_10001) );
oa22f01  g8833 ( .o(n14321), .a(n6966_1), .b(n5705_1), .c(n6959), .d(n14320) );
ao12f01  g8834 ( .o(n14322), .a(n14321), .b(n6585), .c(net_9704) );
ao22f01  g8835 ( .o(n14323), .a(n6582), .b(net_9902), .c(n6577), .d(net_9672) );
ao22f01  g8836 ( .o(n14324), .a(n6590), .b(_net_10033), .c(n6580), .d(net_9803) );
na04f01  g8837 ( .o(n7950), .a(n14324), .b(n14323), .c(n14322), .d(n14319) );
oa12f01  g8838 ( .o(n14326), .a(n7805), .b(n7798), .c(n13886) );
in01f01  g8839 ( .o(n14327), .a(n14326) );
no02f01  g8840 ( .o(n14328), .a(n7809), .b(n7795) );
na02f01  g8841 ( .o(n14329), .a(n14328), .b(n14327) );
in01f01  g8842 ( .o(n14330), .a(n14328) );
na02f01  g8843 ( .o(n14331), .a(n14330), .b(n14326) );
na02f01  g8844 ( .o(n7962), .a(n14331), .b(n14329) );
in01f01  g8845 ( .o(n14333), .a(x3849) );
in01f01  g8846 ( .o(n14334), .a(x3858) );
no02f01  g8847 ( .o(n7967), .a(n14334), .b(n14333) );
oa12f01  g8848 ( .o(n14336), .a(n8865), .b(n13431), .c(n8876_1) );
no02f01  g8849 ( .o(n14337), .a(n8859), .b(n8852) );
in01f01  g8850 ( .o(n14338), .a(n14337) );
na02f01  g8851 ( .o(n14339), .a(n14338), .b(n14336) );
in01f01  g8852 ( .o(n14340), .a(n14336) );
na02f01  g8853 ( .o(n14341), .a(n14337), .b(n14340) );
na02f01  g8854 ( .o(n7972), .a(n14341), .b(n14339) );
no03f01  g8855 ( .o(n14343), .a(n10966), .b(n10964), .c(n10959) );
no02f01  g8856 ( .o(n14344), .a(n10968), .b(n10954) );
in01f01  g8857 ( .o(n14345), .a(n14344) );
ao12f01  g8858 ( .o(n14346), .a(n6746), .b(n14345), .c(n14343) );
oa12f01  g8859 ( .o(n14347), .a(n14346), .b(n14345), .c(n14343) );
na02f01  g8860 ( .o(n14348), .a(n10986), .b(n10967) );
no02f01  g8861 ( .o(n14349), .a(n10987), .b(n10398) );
ao22f01  g8862 ( .o(n14350), .a(n14349), .b(n14348), .c(n6760), .d(_net_10147) );
na02f01  g8863 ( .o(n7977), .a(n14350), .b(n14347) );
ao12f01  g8864 ( .o(n14352), .a(n5658), .b(n6875_1), .c(_net_234) );
ao22f01  g8865 ( .o(n14353), .a(n6878), .b(x5901), .c(n6877), .d(net_9895) );
na02f01  g8866 ( .o(n7982), .a(n14353), .b(n14352) );
na02f01  g8867 ( .o(n14355), .a(n6056), .b(_net_231) );
na02f01  g8868 ( .o(n14356), .a(n6055), .b(net_9959) );
ao22f01  g8869 ( .o(n14357), .a(n6062_1), .b(x6102), .c(n6060), .d(_net_10410) );
na04f01  g8870 ( .o(n7987), .a(n14357), .b(n14356), .c(n14355), .d(n6058) );
ao22f01  g8871 ( .o(n14359), .a(n5842), .b(net_9691), .c(n5841), .d(_net_129) );
na02f01  g8872 ( .o(n14360), .a(n5847), .b(net_9988) );
ao22f01  g8873 ( .o(n14361), .a(n5850), .b(net_9790), .c(n5849_1), .d(net_9889) );
na03f01  g8874 ( .o(n7996), .a(n14361), .b(n14360), .c(n14359) );
na02f01  g8875 ( .o(n14363), .a(n5283), .b(n7991) );
in01f01  g8876 ( .o(n14364), .a(_net_9521) );
no02f01  g8877 ( .o(n14365), .a(n12720), .b(n14364) );
oa12f01  g8878 ( .o(n14366), .a(n7998), .b(n14365), .c(n9462) );
no02f01  g8879 ( .o(n14367), .a(n8002), .b(n14364) );
no02f01  g8880 ( .o(n14368), .a(n14367), .b(n5658) );
na03f01  g8881 ( .o(n8001), .a(n14368), .b(n14366), .c(n14363) );
ao22f01  g8882 ( .o(n14370), .a(n5842), .b(net_9724), .c(n5841), .d(_net_164) );
na02f01  g8883 ( .o(n14371), .a(n5847), .b(net_10021) );
ao22f01  g8884 ( .o(n14372), .a(n5850), .b(net_9823), .c(n5849_1), .d(net_9922) );
na03f01  g8885 ( .o(n8006), .a(n14372), .b(n14371), .c(n14370) );
in01f01  g8886 ( .o(n8011), .a(n7976) );
oa12f01  g8887 ( .o(n8016), .a(n14094), .b(n5498), .c(n5496) );
in01f01  g8888 ( .o(n14376), .a(n7595_1) );
in01f01  g8889 ( .o(n14377), .a(n7588) );
no02f01  g8890 ( .o(n14378), .a(n7589), .b(n14377) );
ao12f01  g8891 ( .o(n14379), .a(n11346), .b(n14378), .c(n14376) );
oa12f01  g8892 ( .o(n14380), .a(n14379), .b(n14378), .c(n14376) );
in01f01  g8893 ( .o(n14381), .a(net_192) );
no02f01  g8894 ( .o(n14382), .a(n14381), .b(_net_191) );
in01f01  g8895 ( .o(n14383), .a(_net_191) );
no02f01  g8896 ( .o(n14384), .a(net_192), .b(n14383) );
oa12f01  g8897 ( .o(n14385), .a(net_9568), .b(n14384), .c(n14382) );
oa12f01  g8898 ( .o(n14386), .a(n14385), .b(n14381), .c(net_9568) );
na02f01  g8899 ( .o(n14387), .a(n11577), .b(n5929) );
in01f01  g8900 ( .o(n14388), .a(n14387) );
ao22f01  g8901 ( .o(n14389), .a(n14388), .b(n14386), .c(n11576), .d(net_101) );
na02f01  g8902 ( .o(n8026), .a(n14389), .b(n14380) );
in01f01  g8903 ( .o(n14391), .a(_net_10201) );
ao12f01  g8904 ( .o(n14392), .a(n5658), .b(n6887), .c(x6028) );
oa12f01  g8905 ( .o(n8031), .a(n14392), .b(n6885_1), .c(n14391) );
in01f01  g8906 ( .o(n14394), .a(net_10292) );
oa22f01  g8907 ( .o(n8036), .a(n9353), .b(n5552_1), .c(n9352), .d(n14394) );
oa22f01  g8908 ( .o(n8041), .a(n7480_1), .b(n5806), .c(n7478), .d(n5546) );
oa22f01  g8909 ( .o(n8046), .a(n5694), .b(n9943), .c(n5692), .d(n5637) );
in01f01  g8910 ( .o(n14398), .a(_net_10322) );
ao12f01  g8911 ( .o(n14399), .a(n5658), .b(n5774), .c(x5003) );
oa12f01  g8912 ( .o(n8051), .a(n14399), .b(n5770), .c(n14398) );
in01f01  g8913 ( .o(n14401), .a(net_10177) );
oa22f01  g8914 ( .o(n8059), .a(n7956), .b(n5567_1), .c(n7955), .d(n14401) );
no02f01  g8915 ( .o(n14403), .a(n8877), .b(n8861) );
in01f01  g8916 ( .o(n14404), .a(n14403) );
oa12f01  g8917 ( .o(n14405), .a(n14404), .b(n8874), .c(n8869) );
na02f01  g8918 ( .o(n14406), .a(n14403), .b(n8875) );
na02f01  g8919 ( .o(n8072), .a(n14406), .b(n14405) );
ao12f01  g8920 ( .o(n14408), .a(n5658), .b(n6875_1), .c(net_243) );
ao22f01  g8921 ( .o(n14409), .a(n6878), .b(x5364), .c(n6877), .d(net_9904) );
na02f01  g8922 ( .o(n8081), .a(n14409), .b(n14408) );
na02f01  g8923 ( .o(n14411), .a(n6025), .b(n7593) );
na02f01  g8924 ( .o(n14412), .a(n14411), .b(n8812) );
oa22f01  g8925 ( .o(n8086), .a(n14412), .b(n8810), .c(n8817), .d(n6025) );
ao12f01  g8926 ( .o(n14414), .a(n5658), .b(n6532), .c(net_253) );
ao22f01  g8927 ( .o(n14415), .a(n6535), .b(x4587), .c(n6534), .d(net_10013) );
na02f01  g8928 ( .o(n8091), .a(n14415), .b(n14414) );
ao22f01  g8929 ( .o(n14417), .a(n11503), .b(x2278), .c(n11502), .d(_net_9405) );
oa12f01  g8930 ( .o(n8096), .a(n14417), .b(n11501), .c(n13101) );
ao12f01  g8931 ( .o(n14419), .a(n5658), .b(n7844), .c(net_248) );
ao22f01  g8932 ( .o(n14420), .a(n7847), .b(x5003), .c(n7846), .d(net_9810) );
na02f01  g8933 ( .o(n8101), .a(n14420), .b(n14419) );
na02f01  g8934 ( .o(n14422), .a(n12761), .b(n7801_1) );
na02f01  g8935 ( .o(n14423), .a(n12762), .b(_net_10119) );
na02f01  g8936 ( .o(n8106), .a(n14423), .b(n14422) );
na02f01  g8937 ( .o(n14425), .a(n7937), .b(net_249) );
na02f01  g8938 ( .o(n14426), .a(n7936), .b(net_9779) );
ao22f01  g8939 ( .o(n14427), .a(n7943), .b(_net_10218), .c(n7942), .d(x4937) );
na04f01  g8940 ( .o(n8111), .a(n14427), .b(n14426), .c(n14425), .d(n7939) );
ao22f01  g8941 ( .o(n14429), .a(n8118), .b(x3071), .c(n8117), .d(_net_9392) );
oa12f01  g8942 ( .o(n8116), .a(n14429), .b(n8116_1), .c(n5696) );
na02f01  g8943 ( .o(n14431), .a(n6056), .b(net_251) );
na02f01  g8944 ( .o(n14432), .a(n6055), .b(net_9979) );
ao22f01  g8945 ( .o(n14433), .a(n6062_1), .b(x4781), .c(n6060), .d(_net_10430) );
na04f01  g8946 ( .o(n8125), .a(n14433), .b(n14432), .c(n14431), .d(n6058) );
in01f01  g8947 ( .o(n14435), .a(_net_10105) );
ao12f01  g8948 ( .o(n14436), .a(n5658), .b(n6160_1), .c(x5498) );
oa12f01  g8949 ( .o(n8130), .a(n14436), .b(n6159), .c(n14435) );
ao12f01  g8950 ( .o(n14438), .a(n8028), .b(n8019), .c(n8021_1) );
no04f01  g8951 ( .o(n14439), .a(n14438), .b(n12589), .c(net_9181), .d(net_9182) );
no02f01  g8952 ( .o(n8135), .a(n14439), .b(n7701) );
na02f01  g8953 ( .o(n14441), .a(n11975), .b(n11378) );
na02f01  g8954 ( .o(n14442), .a(n11976), .b(n11379) );
na03f01  g8955 ( .o(n14443), .a(n14442), .b(n14441), .c(n8638) );
ao12f01  g8956 ( .o(n14444), .a(n7883), .b(n8637), .c(_net_9316) );
na02f01  g8957 ( .o(n8140), .a(n14444), .b(n14443) );
oa12f01  g8958 ( .o(n14446), .a(n6809), .b(n6802), .c(n6798) );
no02f01  g8959 ( .o(n14447), .a(n6812), .b(n6800) );
ao12f01  g8960 ( .o(n14448), .a(n6933), .b(n14447), .c(n14446) );
oa12f01  g8961 ( .o(n14449), .a(n14448), .b(n14447), .c(n14446) );
na02f01  g8962 ( .o(n14450), .a(n6837), .b(n6811_1) );
no02f01  g8963 ( .o(n14451), .a(n6838), .b(n6846_1) );
ao22f01  g8964 ( .o(n14452), .a(n14451), .b(n14450), .c(n6168), .d(_net_10251) );
na02f01  g8965 ( .o(n8145), .a(n14452), .b(n14449) );
na02f01  g8966 ( .o(n14454), .a(n11739), .b(n6937) );
no02f01  g8967 ( .o(n14455), .a(n14454), .b(n11738) );
no03f01  g8968 ( .o(n14456), .a(n14455), .b(n11736), .c(n6163) );
ao22f01  g8969 ( .o(n14457), .a(n6787), .b(_net_10220), .c(n6829), .d(_net_10219) );
no02f01  g8970 ( .o(n14458), .a(n14457), .b(_net_10246) );
ao22f01  g8971 ( .o(n14459), .a(_net_10222), .b(n6780), .c(_net_10221), .d(n6781) );
oa12f01  g8972 ( .o(n14460), .a(n14459), .b(n14457), .c(n8960) );
ao12f01  g8973 ( .o(n14461), .a(n6781), .b(_net_10222), .c(n6780) );
ao22f01  g8974 ( .o(n14462), .a(n14461), .b(n8957), .c(n8969), .d(_net_10248) );
oa12f01  g8975 ( .o(n14463), .a(n14462), .b(n14460), .c(n14458) );
oa22f01  g8976 ( .o(n14464), .a(_net_10251), .b(n9205), .c(n9204), .d(_net_10252) );
in01f01  g8977 ( .o(n14465), .a(n14464) );
ao22f01  g8978 ( .o(n14466), .a(_net_10223), .b(n6807), .c(n6805), .d(_net_10224) );
na03f01  g8979 ( .o(n14467), .a(n14466), .b(n14465), .c(n14463) );
oa22f01  g8980 ( .o(n14468), .a(n9062), .b(n6807), .c(n6828), .d(_net_10223) );
na02f01  g8981 ( .o(n14469), .a(n14468), .b(n14465) );
na03f01  g8982 ( .o(n14470), .a(n14465), .b(_net_10250), .c(n9198) );
ao12f01  g8983 ( .o(n14471), .a(n6811_1), .b(_net_10226), .c(n6813) );
ao22f01  g8984 ( .o(n14472), .a(n14471), .b(n9205), .c(n9204), .d(_net_10252) );
na04f01  g8985 ( .o(n14473), .a(n14472), .b(n14470), .c(n14469), .d(n14467) );
oa22f01  g8986 ( .o(n14474), .a(n9220), .b(_net_10256), .c(_net_10255), .d(n9180) );
oa22f01  g8987 ( .o(n14475), .a(_net_10254), .b(n9172), .c(_net_10253), .d(n8978) );
no02f01  g8988 ( .o(n14476), .a(n14475), .b(n14474) );
na02f01  g8989 ( .o(n14477), .a(n14476), .b(n14473) );
oa12f01  g8990 ( .o(n14478), .a(_net_10253), .b(_net_10254), .c(n9172) );
no03f01  g8991 ( .o(n14479), .a(n14478), .b(n14474), .c(_net_10227) );
no03f01  g8992 ( .o(n14480), .a(n14474), .b(n6770), .c(_net_10228) );
oa12f01  g8993 ( .o(n14481), .a(_net_10255), .b(n9220), .c(_net_10256) );
no02f01  g8994 ( .o(n14482), .a(n14481), .b(_net_10229) );
no03f01  g8995 ( .o(n14483), .a(_net_9851), .b(n6163), .c(n9385) );
oa12f01  g8996 ( .o(n14484), .a(n14483), .b(_net_10230), .c(n6769) );
no04f01  g8997 ( .o(n14485), .a(n14484), .b(n14482), .c(n14480), .d(n14479) );
ao12f01  g8998 ( .o(n14486), .a(n14456), .b(n14485), .c(n14477) );
no04f01  g8999 ( .o(n8150), .a(n14486), .b(_net_10302), .c(net_10304), .d(net_10303) );
na03f01  g9000 ( .o(n14488), .a(n6860), .b(_net_9248), .c(_net_9236) );
oa12f01  g9001 ( .o(n14489), .a(_net_9248), .b(n6500), .c(n6494) );
na03f01  g9002 ( .o(n14490), .a(n6850), .b(n6486), .c(_net_9248) );
ao12f01  g9003 ( .o(n14491), .a(n7852), .b(n10087), .c(n6477) );
ao12f01  g9004 ( .o(n14492), .a(n14491), .b(n6471), .c(_net_9248) );
na04f01  g9005 ( .o(n14493), .a(n14492), .b(n14490), .c(n14489), .d(n14488) );
no02f01  g9006 ( .o(n14494), .a(n6502), .b(n7852) );
ao12f01  g9007 ( .o(n14495), .a(_net_9176), .b(n14494), .c(n6467) );
no02f01  g9008 ( .o(n14496), .a(n14495), .b(n6507_1) );
ao12f01  g9009 ( .o(n14497), .a(_net_9176), .b(n14494), .c(n6483) );
na02f01  g9010 ( .o(n14498), .a(_net_9248), .b(_net_9238) );
oa22f01  g9011 ( .o(n14499), .a(n14498), .b(n6474_1), .c(n14497), .d(n6504) );
no03f01  g9012 ( .o(n14500), .a(n14499), .b(n14496), .c(n14493) );
no02f01  g9013 ( .o(n8155), .a(n14500), .b(n6526_1) );
na02f01  g9014 ( .o(n14502), .a(n6514), .b(net_9618) );
na02f01  g9015 ( .o(n14503), .a(net_313), .b(n6539) );
na04f01  g9016 ( .o(n14504), .a(n14503), .b(n14502), .c(n6541_1), .d(net_9616) );
no02f01  g9017 ( .o(n14505), .a(net_9615), .b(net_313) );
no02f01  g9018 ( .o(n14506), .a(n6542), .b(n6514) );
no02f01  g9019 ( .o(n14507), .a(n14506), .b(n14505) );
no02f01  g9020 ( .o(n14508), .a(n6514), .b(net_9619) );
no02f01  g9021 ( .o(n14509), .a(net_313), .b(n6538) );
no03f01  g9022 ( .o(n14510), .a(net_9620), .b(net_9621), .c(net_9617) );
oa12f01  g9023 ( .o(n14511), .a(n14510), .b(n14509), .c(n14508) );
no03f01  g9024 ( .o(n8160), .a(n14511), .b(n14507), .c(n14504) );
in01f01  g9025 ( .o(n14513), .a(_net_10421) );
ao12f01  g9026 ( .o(n14514), .a(n5658), .b(n6052_1), .c(x5427) );
oa12f01  g9027 ( .o(n8165), .a(n14514), .b(n6048), .c(n14513) );
in01f01  g9028 ( .o(n14516), .a(net_9853) );
oa22f01  g9029 ( .o(n8170), .a(n11258), .b(n10282), .c(n11257), .d(n14516) );
in01f01  g9030 ( .o(n14518), .a(_net_10315) );
ao12f01  g9031 ( .o(n14519), .a(n5658), .b(n5774), .c(x5498) );
oa12f01  g9032 ( .o(n8175), .a(n14519), .b(n5770), .c(n14518) );
in01f01  g9033 ( .o(n14521), .a(net_10087) );
oa22f01  g9034 ( .o(n8180), .a(n6989_1), .b(n5488), .c(n6988), .d(n14521) );
na02f01  g9035 ( .o(n14523), .a(n7742), .b(n7741) );
na03f01  g9036 ( .o(n14524), .a(n14523), .b(n5656), .c(n7744) );
oa12f01  g9037 ( .o(n8185), .a(n14524), .b(n7751), .c(n7742) );
ao12f01  g9038 ( .o(n14526), .a(n5658), .b(n7844), .c(net_237) );
ao22f01  g9039 ( .o(n14527), .a(n7847), .b(x5722), .c(n7846), .d(net_9799) );
na02f01  g9040 ( .o(n8190), .a(n14527), .b(n14526) );
na02f01  g9041 ( .o(n14529), .a(n7358), .b(_net_255) );
na02f01  g9042 ( .o(n14530), .a(n7352), .b(net_9686) );
ao22f01  g9043 ( .o(n14531), .a(n7357), .b(_net_10119), .c(n7353), .d(x4449) );
na04f01  g9044 ( .o(n8195), .a(n14531), .b(n14530), .c(n14529), .d(n7355_1) );
ao22f01  g9045 ( .o(n14533), .a(n11503), .b(x2098), .c(n11502), .d(_net_9408) );
oa12f01  g9046 ( .o(n8200), .a(n14533), .b(n11501), .c(n5696) );
ao22f01  g9047 ( .o(n14535), .a(n11503), .b(x1974), .c(n11502), .d(_net_9410) );
oa12f01  g9048 ( .o(n8205), .a(n14535), .b(n11501), .c(n8114) );
oa22f01  g9049 ( .o(n8214), .a(n7956), .b(n5576), .c(n7955), .d(n6589_1) );
no02f01  g9050 ( .o(n14538), .a(n6724), .b(n6715) );
in01f01  g9051 ( .o(n14539), .a(n14538) );
no02f01  g9052 ( .o(n14540), .a(n14539), .b(n6732) );
na02f01  g9053 ( .o(n14541), .a(n14539), .b(n6732) );
na02f01  g9054 ( .o(n14542), .a(n14541), .b(n10948) );
no02f01  g9055 ( .o(n14543), .a(n6752), .b(_net_10142) );
no03f01  g9056 ( .o(n14544), .a(n14543), .b(n6754), .c(n10398) );
ao12f01  g9057 ( .o(n14545), .a(n14544), .b(n6760), .c(_net_10142) );
oa12f01  g9058 ( .o(n8223), .a(n14545), .b(n14542), .c(n14540) );
na02f01  g9059 ( .o(n14547), .a(n6038), .b(net_241) );
na02f01  g9060 ( .o(n14548), .a(n6037_1), .b(net_9870) );
ao22f01  g9061 ( .o(n14549), .a(n6044), .b(x5498), .c(n6042_1), .d(_net_10315) );
na04f01  g9062 ( .o(n8231), .a(n14549), .b(n14548), .c(n14547), .d(n6040) );
ao12f01  g9063 ( .o(n14551), .a(n5658), .b(n6875_1), .c(net_248) );
ao22f01  g9064 ( .o(n14552), .a(n6878), .b(x5003), .c(n6877), .d(net_9909) );
na02f01  g9065 ( .o(n8240), .a(n14552), .b(n14551) );
oa22f01  g9066 ( .o(n8245), .a(n5694), .b(n5821), .c(n5692), .d(n5546) );
oa22f01  g9067 ( .o(n8250), .a(n5907), .b(n9009), .c(n5905), .d(n5637) );
in01f01  g9068 ( .o(n14556), .a(net_10186) );
oa22f01  g9069 ( .o(n8255), .a(n7956), .b(n5640), .c(n7955), .d(n14556) );
no02f01  g9070 ( .o(n14558), .a(n9186), .b(n9177) );
na02f01  g9071 ( .o(n14559), .a(n14558), .b(n9214) );
in01f01  g9072 ( .o(n14560), .a(n14558) );
oa12f01  g9073 ( .o(n14561), .a(n14560), .b(n9213), .c(n9211) );
na02f01  g9074 ( .o(n8260), .a(n14561), .b(n14559) );
in01f01  g9075 ( .o(n14563), .a(n8966) );
no02f01  g9076 ( .o(n14564), .a(n8959), .b(n8958) );
in01f01  g9077 ( .o(n14565), .a(n14564) );
na02f01  g9078 ( .o(n14566), .a(n14565), .b(n14563) );
na02f01  g9079 ( .o(n14567), .a(n14564), .b(n8966) );
na02f01  g9080 ( .o(n8268), .a(n14567), .b(n14566) );
in01f01  g9081 ( .o(n14569), .a(net_10395) );
oa22f01  g9082 ( .o(n8276), .a(n10211), .b(n5546), .c(n10210), .d(n14569) );
ao12f01  g9083 ( .o(n14571), .a(n5658), .b(n6532), .c(net_257) );
ao22f01  g9084 ( .o(n14572), .a(n6535), .b(x4285), .c(n6534), .d(net_10017) );
na02f01  g9085 ( .o(n8281), .a(n14572), .b(n14571) );
na02f01  g9086 ( .o(n14574), .a(n12555), .b(net_9277) );
na02f01  g9087 ( .o(n14575), .a(n12554), .b(n12550) );
ao12f01  g9088 ( .o(n8286), .a(n10005), .b(n14575), .c(n14574) );
in01f01  g9089 ( .o(n14577), .a(_net_10213) );
ao12f01  g9090 ( .o(n14578), .a(n5658), .b(n6887), .c(x5289) );
oa12f01  g9091 ( .o(n8291), .a(n14578), .b(n6885_1), .c(n14577) );
ao12f01  g9092 ( .o(n14580), .a(n5658), .b(n6532), .c(net_239) );
ao22f01  g9093 ( .o(n14581), .a(n6535), .b(x5601), .c(n6534), .d(net_9999) );
na02f01  g9094 ( .o(n8296), .a(n14581), .b(n14580) );
no02f01  g9095 ( .o(n8301), .a(n11346), .b(n6009_1) );
oa22f01  g9096 ( .o(n8310), .a(n11882), .b(n8686), .c(n11881), .d(n12510) );
na02f01  g9097 ( .o(n14585), .a(n8091_1), .b(n8547) );
na02f01  g9098 ( .o(n14586), .a(n14585), .b(n9399) );
oa22f01  g9099 ( .o(n8315), .a(n14586), .b(n9397), .c(n9407), .d(n8091_1) );
na02f01  g9100 ( .o(n14588), .a(n7937), .b(net_240) );
na02f01  g9101 ( .o(n14589), .a(n7936), .b(net_9770) );
ao22f01  g9102 ( .o(n14590), .a(n7943), .b(_net_10209), .c(n7942), .d(x5548) );
na04f01  g9103 ( .o(n8320), .a(n14590), .b(n14589), .c(n14588), .d(n7939) );
na02f01  g9104 ( .o(n14592), .a(n6038), .b(_net_234) );
na02f01  g9105 ( .o(n14593), .a(n6037_1), .b(net_9863) );
ao22f01  g9106 ( .o(n14594), .a(n6044), .b(x5901), .c(n6042_1), .d(_net_10308) );
na04f01  g9107 ( .o(n8325), .a(n14594), .b(n14593), .c(n14592), .d(n6040) );
oa22f01  g9108 ( .o(n8330), .a(n7738_1), .b(n6454), .c(n7736), .d(n8339_1) );
in01f01  g9109 ( .o(n14597), .a(net_10187) );
oa22f01  g9110 ( .o(n8335), .a(n7956), .b(n5552_1), .c(n7955), .d(n14597) );
na02f01  g9111 ( .o(n14599), .a(n7670_1), .b(_net_10435) );
na02f01  g9112 ( .o(n8344), .a(n14599), .b(n7672) );
oa22f01  g9113 ( .o(n8349), .a(n7367), .b(n6596), .c(n7365_1), .d(n5576) );
ao22f01  g9114 ( .o(n14602), .a(n5842), .b(net_9674), .c(n5841), .d(net_112) );
na02f01  g9115 ( .o(n14603), .a(n5847), .b(net_9971) );
ao22f01  g9116 ( .o(n14604), .a(n5850), .b(net_9773), .c(n5849_1), .d(net_9872) );
na03f01  g9117 ( .o(n8354), .a(n14604), .b(n14603), .c(n14602) );
ao12f01  g9118 ( .o(n14606), .a(n5658), .b(n5678), .c(net_257) );
ao22f01  g9119 ( .o(n14607), .a(n5681_1), .b(x4285), .c(n5680), .d(net_9720) );
na02f01  g9120 ( .o(n8358), .a(n14607), .b(n14606) );
na03f01  g9121 ( .o(n14609), .a(_net_10221), .b(_net_10220), .c(_net_10219) );
na02f01  g9122 ( .o(n8363), .a(n14609), .b(n9064) );
in01f01  g9123 ( .o(n14611), .a(_net_10214) );
ao12f01  g9124 ( .o(n14612), .a(n5658), .b(n6887), .c(x5225) );
oa12f01  g9125 ( .o(n8372), .a(n14612), .b(n6885_1), .c(n14611) );
no02f01  g9126 ( .o(n14614), .a(n8904), .b(n8888) );
in01f01  g9127 ( .o(n14615), .a(n14614) );
na02f01  g9128 ( .o(n14616), .a(n14615), .b(n10676) );
na03f01  g9129 ( .o(n14617), .a(n14614), .b(n8881), .c(n8856) );
na02f01  g9130 ( .o(n8384), .a(n14617), .b(n14616) );
oa22f01  g9131 ( .o(n8389), .a(n7756), .b(n5791), .c(n7755), .d(n12262) );
na02f01  g9132 ( .o(n14620), .a(n6175), .b(n6172) );
na02f01  g9133 ( .o(n14621), .a(n6172), .b(n6183) );
na03f01  g9134 ( .o(n14622), .a(n14621), .b(n6186_1), .c(n6177_1) );
na02f01  g9135 ( .o(n14623), .a(n6168), .b(_net_10257) );
na03f01  g9136 ( .o(n8394), .a(n14623), .b(n14622), .c(n14620) );
ao22f01  g9137 ( .o(n14625), .a(_net_10233), .b(n6781), .c(_net_10234), .d(n6780) );
no02f01  g9138 ( .o(n14626), .a(_net_10232), .b(n6787) );
ao22f01  g9139 ( .o(n14627), .a(_net_10232), .b(n6787), .c(n6829), .d(_net_8843) );
oa12f01  g9140 ( .o(n14628), .a(n14625), .b(n14627), .c(n14626) );
in01f01  g9141 ( .o(n14629), .a(_net_10234) );
in01f01  g9142 ( .o(n14630), .a(_net_10233) );
ao12f01  g9143 ( .o(n14631), .a(n6781), .b(_net_10234), .c(n6780) );
ao22f01  g9144 ( .o(n14632), .a(n14631), .b(n14630), .c(n14629), .d(_net_10248) );
ao22f01  g9145 ( .o(n14633), .a(n6811_1), .b(net_10237), .c(net_10238), .d(n6813) );
ao22f01  g9146 ( .o(n14634), .a(_net_10236), .b(n6805), .c(_net_10235), .d(n6807) );
na02f01  g9147 ( .o(n14635), .a(n14634), .b(n14633) );
ao12f01  g9148 ( .o(n14636), .a(n14635), .b(n14632), .c(n14628) );
in01f01  g9149 ( .o(n14637), .a(net_10240) );
oa12f01  g9150 ( .o(n14638), .a(_net_10253), .b(_net_10254), .c(n14637) );
oa22f01  g9151 ( .o(n14639), .a(n14638), .b(net_10239), .c(n6770), .d(net_10240) );
ao22f01  g9152 ( .o(n14640), .a(_net_10241), .b(n11506), .c(_net_10242), .d(n6769) );
in01f01  g9153 ( .o(n14641), .a(_net_10242) );
oa12f01  g9154 ( .o(n14642), .a(_net_10255), .b(n14641), .c(_net_10256) );
oa22f01  g9155 ( .o(n14643), .a(n14642), .b(_net_10241), .c(_net_10242), .d(n6769) );
ao12f01  g9156 ( .o(n14644), .a(n14643), .b(n14640), .c(n14639) );
in01f01  g9157 ( .o(n14645), .a(_net_10236) );
oa12f01  g9158 ( .o(n14646), .a(_net_10249), .b(n14645), .c(_net_10250) );
oa22f01  g9159 ( .o(n14647), .a(n14646), .b(_net_10235), .c(_net_10236), .d(n6805) );
in01f01  g9160 ( .o(n14648), .a(net_10238) );
oa12f01  g9161 ( .o(n14649), .a(_net_10251), .b(n14648), .c(_net_10252) );
oa22f01  g9162 ( .o(n14650), .a(n14649), .b(net_10237), .c(net_10238), .d(n6813) );
ao12f01  g9163 ( .o(n14651), .a(n14650), .b(n14647), .c(n14633) );
na02f01  g9164 ( .o(n14652), .a(n14651), .b(n14644) );
in01f01  g9165 ( .o(n14653), .a(n14640) );
in01f01  g9166 ( .o(n14654), .a(net_10239) );
oa22f01  g9167 ( .o(n14655), .a(_net_10254), .b(n14637), .c(_net_10253), .d(n14654) );
oa12f01  g9168 ( .o(n14656), .a(n14644), .b(n14655), .c(n14653) );
oa12f01  g9169 ( .o(n8399), .a(n14656), .b(n14652), .c(n14636) );
no02f01  g9170 ( .o(n14658), .a(n12420), .b(n12404) );
no02f01  g9171 ( .o(n14659), .a(n12402), .b(n12401) );
na02f01  g9172 ( .o(n14660), .a(n14659), .b(n14658) );
in01f01  g9173 ( .o(n14661), .a(n14659) );
oa12f01  g9174 ( .o(n14662), .a(n14661), .b(n12420), .c(n12404) );
na02f01  g9175 ( .o(n8404), .a(n14662), .b(n14660) );
na02f01  g9176 ( .o(n14664), .a(n11860), .b(n8087) );
na02f01  g9177 ( .o(n14665), .a(n11859), .b(_net_9217) );
na02f01  g9178 ( .o(n14666), .a(n14665), .b(n14664) );
oa22f01  g9179 ( .o(n8409), .a(n14666), .b(n9397), .c(n9407), .d(n8087) );
oa22f01  g9180 ( .o(n8414), .a(n8418), .b(n8725), .c(n8417), .d(n5570) );
ao12f01  g9181 ( .o(n14669), .a(n5658), .b(n7844), .c(net_235) );
ao22f01  g9182 ( .o(n14670), .a(n7847), .b(x5850), .c(n7846), .d(net_9797) );
na02f01  g9183 ( .o(n8419), .a(n14670), .b(n14669) );
ao22f01  g9184 ( .o(n14672), .a(n5842), .b(net_9713), .c(n5841), .d(_net_153) );
na02f01  g9185 ( .o(n14673), .a(n5847), .b(net_10010) );
ao22f01  g9186 ( .o(n14674), .a(n5850), .b(net_9812), .c(n5849_1), .d(net_9911) );
na03f01  g9187 ( .o(n8424), .a(n14674), .b(n14673), .c(n14672) );
no02f01  g9188 ( .o(n8429), .a(n9566), .b(n5927) );
na02f01  g9189 ( .o(n14677), .a(n6349), .b(n6265) );
oa22f01  g9190 ( .o(n8438), .a(n14677), .b(n6348), .c(n6349), .d(n8870) );
no02f01  g9191 ( .o(n14679), .a(n7305), .b(n7234) );
no02f01  g9192 ( .o(n14680), .a(n7274), .b(n7203) );
no02f01  g9193 ( .o(n14681), .a(n14680), .b(n14679) );
no02f01  g9194 ( .o(n14682), .a(n14681), .b(n10248) );
na02f01  g9195 ( .o(n14683), .a(n14681), .b(n10248) );
na02f01  g9196 ( .o(n14684), .a(n14683), .b(n6148) );
ao12f01  g9197 ( .o(n14685), .a(n6131_1), .b(n6147), .c(net_9366) );
oa12f01  g9198 ( .o(n8447), .a(n14685), .b(n14684), .c(n14682) );
na02f01  g9199 ( .o(n14687), .a(n7425), .b(n7370_1) );
na03f01  g9200 ( .o(n14688), .a(n14687), .b(n7431), .c(n7427) );
oa12f01  g9201 ( .o(n14689), .a(n7450), .b(n7446_1), .c(_net_10477) );
ao12f01  g9202 ( .o(n14690), .a(n14689), .b(n7446_1), .c(_net_10477) );
ao12f01  g9203 ( .o(n14691), .a(n14690), .b(n7453), .c(_net_10477) );
na02f01  g9204 ( .o(n8452), .a(n14691), .b(n14688) );
in01f01  g9205 ( .o(n14693), .a(net_10388) );
oa22f01  g9206 ( .o(n8457), .a(n10211), .b(n5609), .c(n10210), .d(n14693) );
oa12f01  g9207 ( .o(n14695), .a(n8912), .b(n13995), .c(_net_9600) );
in01f01  g9208 ( .o(n14696), .a(n14695) );
ao12f01  g9209 ( .o(n14697), .a(n14696), .b(n13995), .c(_net_9600) );
no03f01  g9210 ( .o(n14698), .a(n13998), .b(n13991), .c(n6653) );
in01f01  g9211 ( .o(n14699), .a(_net_9601) );
no02f01  g9212 ( .o(n14700), .a(n8918), .b(n14699) );
no02f01  g9213 ( .o(n14701), .a(n6014), .b(_net_9601) );
no02f01  g9214 ( .o(n14702), .a(n14701), .b(n14700) );
oa12f01  g9215 ( .o(n14703), .a(n14702), .b(n14698), .c(n14697) );
no02f01  g9216 ( .o(n14704), .a(n14698), .b(n14697) );
in01f01  g9217 ( .o(n14705), .a(n14702) );
na02f01  g9218 ( .o(n14706), .a(n14705), .b(n14704) );
na02f01  g9219 ( .o(n8462), .a(n14706), .b(n14703) );
ao22f01  g9220 ( .o(n14708), .a(n5842), .b(net_9690), .c(n5841), .d(_net_128) );
na02f01  g9221 ( .o(n14709), .a(n5847), .b(net_9987) );
ao22f01  g9222 ( .o(n14710), .a(n5850), .b(net_9789), .c(n5849_1), .d(net_9888) );
na03f01  g9223 ( .o(n8467), .a(n14710), .b(n14709), .c(n14708) );
in01f01  g9224 ( .o(n14712), .a(x3683) );
in01f01  g9225 ( .o(n14713), .a(net_9162) );
na04f01  g9226 ( .o(n14714), .a(_net_9118), .b(n14713), .c(n14712), .d(x6599) );
na03f01  g9227 ( .o(n14715), .a(n14713), .b(x3683), .c(x6599) );
na02f01  g9228 ( .o(n8472), .a(n14715), .b(n14714) );
no02f01  g9229 ( .o(n14717), .a(n10390), .b(_net_10162) );
na02f01  g9230 ( .o(n14718), .a(n10391), .b(n10948) );
oa12f01  g9231 ( .o(n14719), .a(n6750), .b(n10396), .c(_net_10162) );
ao12f01  g9232 ( .o(n14720), .a(n14719), .b(n10396), .c(_net_10162) );
ao12f01  g9233 ( .o(n14721), .a(n14720), .b(n6760), .c(_net_10162) );
oa12f01  g9234 ( .o(n8477), .a(n14721), .b(n14718), .c(n14717) );
na03f01  g9235 ( .o(n14723), .a(n10045), .b(n6130), .c(_net_9382) );
na03f01  g9236 ( .o(n14724), .a(n10894), .b(n6140), .c(_net_9382) );
na03f01  g9237 ( .o(n14725), .a(n10897), .b(_net_9382), .c(n6136_1) );
na02f01  g9238 ( .o(n14726), .a(n8105), .b(n6136_1) );
ao12f01  g9239 ( .o(n14727), .a(n5658), .b(n14726), .c(_net_9385) );
na04f01  g9240 ( .o(n8482), .a(n14727), .b(n14725), .c(n14724), .d(n14723) );
no03f01  g9241 ( .o(n14729), .a(n7594), .b(n7591), .c(net_9545) );
na02f01  g9242 ( .o(n14730), .a(n11345), .b(n7595_1) );
no02f01  g9243 ( .o(n14731), .a(net_9568), .b(_net_191) );
no02f01  g9244 ( .o(n14732), .a(n8578), .b(n14383) );
no02f01  g9245 ( .o(n14733), .a(n14732), .b(n14731) );
ao22f01  g9246 ( .o(n14734), .a(n14733), .b(n14388), .c(n11576), .d(net_100) );
oa12f01  g9247 ( .o(n8491), .a(n14734), .b(n14730), .c(n14729) );
ao12f01  g9248 ( .o(n14736), .a(n5658), .b(n6532), .c(net_246) );
ao22f01  g9249 ( .o(n14737), .a(n6535), .b(x5143), .c(n6534), .d(net_10006) );
na02f01  g9250 ( .o(n8496), .a(n14737), .b(n14736) );
in01f01  g9251 ( .o(n14739), .a(n8899) );
in01f01  g9252 ( .o(n14740), .a(n8884) );
oa12f01  g9253 ( .o(n14741), .a(n14740), .b(n12748), .c(n8907) );
na02f01  g9254 ( .o(n14742), .a(n14741), .b(n14739) );
no02f01  g9255 ( .o(n14743), .a(n8900), .b(n8883) );
in01f01  g9256 ( .o(n14744), .a(n14743) );
na02f01  g9257 ( .o(n14745), .a(n14744), .b(n14742) );
na03f01  g9258 ( .o(n14746), .a(n14743), .b(n14741), .c(n14739) );
na02f01  g9259 ( .o(n8505), .a(n14746), .b(n14745) );
in01f01  g9260 ( .o(n14748), .a(_net_165) );
oa12f01  g9261 ( .o(n8510), .a(n14748), .b(n11920), .c(n11916) );
ao22f01  g9262 ( .o(n14750), .a(n5842), .b(net_9670), .c(n5841), .d(net_108) );
na02f01  g9263 ( .o(n14751), .a(n5847), .b(net_9967) );
ao22f01  g9264 ( .o(n14752), .a(n5850), .b(net_9769), .c(n5849_1), .d(net_9868) );
na03f01  g9265 ( .o(n8515), .a(n14752), .b(n14751), .c(n14750) );
no02f01  g9266 ( .o(n14754), .a(n8705), .b(net_9655) );
no03f01  g9267 ( .o(n8519), .a(n14754), .b(n10525), .c(net_9151) );
in01f01  g9268 ( .o(n14756), .a(_net_10211) );
ao12f01  g9269 ( .o(n14757), .a(n5658), .b(n6887), .c(x5427) );
oa12f01  g9270 ( .o(n8524), .a(n14757), .b(n6885_1), .c(n14756) );
ao22f01  g9271 ( .o(n14759), .a(n6602), .b(net_10006), .c(n6597), .d(_net_9740) );
ao22f01  g9272 ( .o(n14760), .a(n6577), .b(net_9677), .c(n6555), .d(net_9974) );
in01f01  g9273 ( .o(n14761), .a(net_9808) );
oa22f01  g9274 ( .o(n14762), .a(n6966_1), .b(n8181), .c(n9978), .d(n14761) );
na02f01  g9275 ( .o(n14763), .a(n6585), .b(net_9709) );
na02f01  g9276 ( .o(n14764), .a(n6582), .b(net_9907) );
na02f01  g9277 ( .o(n14765), .a(n14764), .b(n14763) );
ao22f01  g9278 ( .o(n14766), .a(n6590), .b(_net_10037), .c(n6573), .d(net_9875) );
ao22f01  g9279 ( .o(n14767), .a(n6599_1), .b(_net_9839), .c(n6584_1), .d(net_9776) );
na02f01  g9280 ( .o(n14768), .a(n14767), .b(n14766) );
no03f01  g9281 ( .o(n14769), .a(n14768), .b(n14765), .c(n14762) );
na03f01  g9282 ( .o(n8534), .a(n14769), .b(n14760), .c(n14759) );
ao12f01  g9283 ( .o(n14771), .a(n5658), .b(n7844), .c(net_238) );
ao22f01  g9284 ( .o(n14772), .a(n7847), .b(x5647), .c(n7846), .d(net_9800) );
na02f01  g9285 ( .o(n8538), .a(n14772), .b(n14771) );
oa22f01  g9286 ( .o(n8543), .a(n5907), .b(n7389_1), .c(n5905), .d(n5573) );
no02f01  g9287 ( .o(n14775), .a(n13122), .b(n5658) );
oa12f01  g9288 ( .o(n14776), .a(n14775), .b(n5693), .c(x4587) );
oa12f01  g9289 ( .o(n8548), .a(n14776), .b(n13123), .c(n13776) );
ao22f01  g9290 ( .o(n14778), .a(n5842), .b(net_9727), .c(n5841), .d(_net_168) );
na02f01  g9291 ( .o(n14779), .a(n5847), .b(net_10024) );
ao22f01  g9292 ( .o(n14780), .a(n5850), .b(net_9826), .c(n5849_1), .d(net_9925) );
na03f01  g9293 ( .o(n8553), .a(n14780), .b(n14779), .c(n14778) );
ao22f01  g9294 ( .o(n14782), .a(n5842), .b(_net_9728), .c(n5841), .d(_net_169) );
na02f01  g9295 ( .o(n14783), .a(n5847), .b(_net_10025) );
ao22f01  g9296 ( .o(n14784), .a(n5850), .b(_net_9827), .c(n5849_1), .d(_net_9926) );
na03f01  g9297 ( .o(n8558), .a(n14784), .b(n14783), .c(n14782) );
na02f01  g9298 ( .o(n14786), .a(n5935_1), .b(_net_9567) );
ao12f01  g9299 ( .o(n14787), .a(_net_9565), .b(n6009_1), .c(net_9570) );
na02f01  g9300 ( .o(n8567), .a(n14787), .b(n14786) );
no02f01  g9301 ( .o(n14789), .a(n9910), .b(net_9221) );
no03f01  g9302 ( .o(n8572), .a(n14789), .b(n9912), .c(n9904) );
in01f01  g9303 ( .o(n14791), .a(net_9620) );
no03f01  g9304 ( .o(n14792), .a(n6548), .b(n14791), .c(n6538) );
oa12f01  g9305 ( .o(n14793), .a(n6550), .b(n14792), .c(net_9621) );
ao12f01  g9306 ( .o(n8582), .a(n14793), .b(n14792), .c(net_9621) );
in01f01  g9307 ( .o(n14795), .a(_net_10091) );
ao12f01  g9308 ( .o(n8587), .a(n6155_1), .b(n10699), .c(n14795) );
oa22f01  g9309 ( .o(n8592), .a(n7480_1), .b(n6904), .c(n7478), .d(n5537_1) );
na02f01  g9310 ( .o(n14798), .a(_net_10220), .b(n3465) );
na02f01  g9311 ( .o(n14799), .a(n8960), .b(_net_10219) );
na02f01  g9312 ( .o(n8597), .a(n14799), .b(n14798) );
no02f01  g9313 ( .o(n14801), .a(n6549), .b(net_9620) );
no03f01  g9314 ( .o(n8602), .a(n14801), .b(n14792), .c(net_9613) );
ao12f01  g9315 ( .o(n14803), .a(n5658), .b(n6532), .c(_net_232) );
ao22f01  g9316 ( .o(n14804), .a(n6535), .b(x6028), .c(n6534), .d(net_9992) );
na02f01  g9317 ( .o(n8607), .a(n14804), .b(n14803) );
ao22f01  g9318 ( .o(n14806), .a(n5842), .b(net_9696), .c(n5841), .d(net_136) );
na02f01  g9319 ( .o(n14807), .a(n5847), .b(net_9993) );
ao22f01  g9320 ( .o(n14808), .a(n5850), .b(net_9795), .c(n5849_1), .d(net_9894) );
na03f01  g9321 ( .o(n8612), .a(n14808), .b(n14807), .c(n14806) );
in01f01  g9322 ( .o(n14810), .a(net_225) );
oa22f01  g9323 ( .o(n8616), .a(n8418), .b(n14810), .c(n8417), .d(n5513_1) );
na02f01  g9324 ( .o(n14812), .a(n6349), .b(n6305) );
oa22f01  g9325 ( .o(n8626), .a(n14812), .b(n6348), .c(n6349), .d(n8898) );
ao12f01  g9326 ( .o(n14814), .a(n5658), .b(n6052_1), .c(x4587) );
oa12f01  g9327 ( .o(n8631), .a(n14814), .b(n6048), .c(n8219_1) );
no02f01  g9328 ( .o(n14816), .a(n9551), .b(n8756) );
na03f01  g9329 ( .o(n14817), .a(n14816), .b(_net_9611), .c(_net_9641) );
no02f01  g9330 ( .o(n8636), .a(n14817), .b(n9490) );
na02f01  g9331 ( .o(n14819), .a(n6836), .b(n7991) );
na02f01  g9332 ( .o(n14820), .a(_net_9517), .b(_net_9516) );
ao12f01  g9333 ( .o(n14821), .a(n7999), .b(n14820), .c(n7987_1) );
in01f01  g9334 ( .o(n14822), .a(_net_9517) );
oa12f01  g9335 ( .o(n14823), .a(x6599), .b(n8002), .c(n14822) );
no02f01  g9336 ( .o(n14824), .a(n14823), .b(n14821) );
na02f01  g9337 ( .o(n8641), .a(n14824), .b(n14819) );
ao12f01  g9338 ( .o(n14826), .a(n5658), .b(n6887), .c(x4587) );
oa12f01  g9339 ( .o(n8650), .a(n14826), .b(n6885_1), .c(n8969) );
oa22f01  g9340 ( .o(n14828), .a(n13697), .b(n10693), .c(n10694), .d(n11492) );
ao12f01  g9341 ( .o(n14829), .a(n14828), .b(net_10078), .c(net_10069) );
oa22f01  g9342 ( .o(n14830), .a(n10699), .b(n10520), .c(n10462), .d(n8667) );
oa22f01  g9343 ( .o(n14831), .a(n13973), .b(n10701), .c(n13732), .d(n6152) );
no02f01  g9344 ( .o(n14832), .a(n14831), .b(n14830) );
no04f01  g9345 ( .o(n14833), .a(_net_9957), .b(_net_10056), .c(net_9858), .d(net_9759) );
ao22f01  g9346 ( .o(n14834), .a(net_10071), .b(net_10080), .c(net_10063), .d(net_10072) );
na04f01  g9347 ( .o(n8655), .a(n14834), .b(n14833), .c(n14832), .d(n14829) );
na02f01  g9348 ( .o(n14836), .a(n6056), .b(_net_255) );
na02f01  g9349 ( .o(n14837), .a(n6055), .b(net_9983) );
ao22f01  g9350 ( .o(n14838), .a(n6062_1), .b(x4449), .c(n6060), .d(_net_10434) );
na04f01  g9351 ( .o(n8659), .a(n14838), .b(n14837), .c(n14836), .d(n6058) );
ao22f01  g9352 ( .o(n14840), .a(n8047), .b(net_10064), .c(n6564), .d(net_10086) );
oa12f01  g9353 ( .o(n14841), .a(n14840), .b(n6563), .c(n9518) );
in01f01  g9354 ( .o(n14842), .a(net_9814) );
oa22f01  g9355 ( .o(n14843), .a(n6593), .b(n14597), .c(n9978), .d(n14842) );
oa22f01  g9356 ( .o(n14844), .a(n8302), .b(n14394), .c(n6600), .d(n5797_1) );
no03f01  g9357 ( .o(n14845), .a(n14844), .b(n14843), .c(n14841) );
ao22f01  g9358 ( .o(n14846), .a(n6606), .b(_net_9944), .c(n6597), .d(_net_9746) );
ao22f01  g9359 ( .o(n14847), .a(n6585), .b(net_9715), .c(n6584_1), .d(net_9782) );
na02f01  g9360 ( .o(n14848), .a(n6582), .b(net_9913) );
na02f01  g9361 ( .o(n14849), .a(n6602), .b(net_10012) );
na02f01  g9362 ( .o(n14850), .a(n14849), .b(n14848) );
na02f01  g9363 ( .o(n14851), .a(n6573), .b(net_9881) );
oa12f01  g9364 ( .o(n14852), .a(n14851), .b(n6591), .c(n5827) );
in01f01  g9365 ( .o(n14853), .a(net_9980) );
oa22f01  g9366 ( .o(n14854), .a(n11677), .b(n12055), .c(n6955), .d(n14853) );
na02f01  g9367 ( .o(n14855), .a(n6577), .b(net_9683) );
oa12f01  g9368 ( .o(n14856), .a(n14855), .b(n8299), .c(n7463) );
no04f01  g9369 ( .o(n14857), .a(n14856), .b(n14854), .c(n14852), .d(n14850) );
na04f01  g9370 ( .o(n8664), .a(n14857), .b(n14847), .c(n14846), .d(n14845) );
in01f01  g9371 ( .o(n14859), .a(n7980) );
na02f01  g9372 ( .o(n14860), .a(n14822), .b(_net_9516) );
no04f01  g9373 ( .o(n14861), .a(n14860), .b(n7985), .c(n7983), .d(n5877) );
na04f01  g9374 ( .o(n14862), .a(n7989), .b(n14859), .c(_net_9514), .d(x6599) );
oa22f01  g9375 ( .o(n8668), .a(n14862), .b(n14861), .c(n14859), .d(n5658) );
na02f01  g9376 ( .o(n14864), .a(n9948), .b(n8189) );
no02f01  g9377 ( .o(n14865), .a(n14864), .b(n9947) );
no03f01  g9378 ( .o(n14866), .a(n14865), .b(n9945), .c(n8181) );
ao22f01  g9379 ( .o(n14867), .a(_net_10325), .b(n9128), .c(n9129), .d(_net_10324) );
no02f01  g9380 ( .o(n14868), .a(n14867), .b(_net_10351) );
ao22f01  g9381 ( .o(n14869), .a(n9089), .b(_net_10327), .c(n9087), .d(_net_10326) );
oa12f01  g9382 ( .o(n14870), .a(n14869), .b(n14867), .c(n7027) );
ao12f01  g9383 ( .o(n14871), .a(n9087), .b(n9089), .c(_net_10327) );
ao22f01  g9384 ( .o(n14872), .a(n14871), .b(n7018), .c(_net_10353), .d(n7017_1) );
oa12f01  g9385 ( .o(n14873), .a(n14872), .b(n14870), .c(n14868) );
oa22f01  g9386 ( .o(n14874), .a(_net_10356), .b(n7049), .c(_net_10357), .d(n7048_1) );
in01f01  g9387 ( .o(n14875), .a(n14874) );
ao22f01  g9388 ( .o(n14876), .a(_net_10329), .b(n9104), .c(n9106), .d(_net_10328) );
na03f01  g9389 ( .o(n14877), .a(n14876), .b(n14875), .c(n14873) );
oa22f01  g9390 ( .o(n14878), .a(n9127), .b(_net_10328), .c(n8933), .d(n9106) );
na02f01  g9391 ( .o(n14879), .a(n14878), .b(n14875) );
na03f01  g9392 ( .o(n14880), .a(n14875), .b(n7042), .c(_net_10355) );
ao12f01  g9393 ( .o(n14881), .a(n9110), .b(n9112), .c(_net_10331) );
ao22f01  g9394 ( .o(n14882), .a(n14881), .b(n7049), .c(_net_10357), .d(n7048_1) );
na04f01  g9395 ( .o(n14883), .a(n14882), .b(n14880), .c(n14879), .d(n14877) );
oa22f01  g9396 ( .o(n14884), .a(_net_10360), .b(n7064), .c(n8931), .d(_net_10361) );
oa22f01  g9397 ( .o(n14885), .a(n6999), .b(_net_10358), .c(n6994), .d(_net_10359) );
no02f01  g9398 ( .o(n14886), .a(n14885), .b(n14884) );
na02f01  g9399 ( .o(n14887), .a(n14886), .b(n14883) );
oa12f01  g9400 ( .o(n14888), .a(_net_10358), .b(n6994), .c(_net_10359) );
no03f01  g9401 ( .o(n14889), .a(n14888), .b(n14884), .c(_net_10332) );
no03f01  g9402 ( .o(n14890), .a(n14884), .b(_net_10333), .c(n9077) );
oa12f01  g9403 ( .o(n14891), .a(_net_10360), .b(n8931), .c(_net_10361) );
no02f01  g9404 ( .o(n14892), .a(n14891), .b(_net_10334) );
no03f01  g9405 ( .o(n14893), .a(_net_9950), .b(n9579), .c(n8181) );
oa12f01  g9406 ( .o(n14894), .a(n14893), .b(_net_10335), .c(n10140) );
no04f01  g9407 ( .o(n14895), .a(n14894), .b(n14892), .c(n14890), .d(n14889) );
ao12f01  g9408 ( .o(n14896), .a(n14866), .b(n14895), .c(n14887) );
no04f01  g9409 ( .o(n8673), .a(n14896), .b(_net_10407), .c(net_10408), .d(net_10409) );
ao12f01  g9410 ( .o(n14898), .a(n5658), .b(n6532), .c(net_235) );
ao22f01  g9411 ( .o(n14899), .a(n6535), .b(x5850), .c(n6534), .d(net_9995) );
na02f01  g9412 ( .o(n8678), .a(n14899), .b(n14898) );
oa22f01  g9413 ( .o(n8683), .a(n7480_1), .b(n8583), .c(n7478), .d(n5570) );
no03f01  g9414 ( .o(n14902), .a(n6517_1), .b(n6513), .c(n8509) );
no02f01  g9415 ( .o(n14903), .a(n14902), .b(n6673) );
no02f01  g9416 ( .o(n14904), .a(n14903), .b(n6511) );
in01f01  g9417 ( .o(n14905), .a(n6472) );
na03f01  g9418 ( .o(n14906), .a(n6467), .b(n6464_1), .c(_net_9244) );
ao12f01  g9419 ( .o(n14907), .a(n6463), .b(n14906), .c(n14905) );
na02f01  g9420 ( .o(n14908), .a(n6471), .b(_net_9244) );
oa12f01  g9421 ( .o(n14909), .a(_net_9244), .b(n10086), .c(n6476) );
oa12f01  g9422 ( .o(n14910), .a(n14909), .b(n14908), .c(n7852) );
no03f01  g9423 ( .o(n14911), .a(n14910), .b(n14907), .c(n14904) );
oa12f01  g9424 ( .o(n14912), .a(_net_9244), .b(n6483), .c(n6480) );
ao12f01  g9425 ( .o(n14913), .a(n6479_1), .b(n14912), .c(n6486) );
ao12f01  g9426 ( .o(n14914), .a(n8509), .b(n6499), .c(n6493_1) );
ao12f01  g9427 ( .o(n14915), .a(n14908), .b(n7863), .c(n7862_1) );
no03f01  g9428 ( .o(n14916), .a(n14915), .b(n14914), .c(n14913) );
ao12f01  g9429 ( .o(n8688), .a(n6526_1), .b(n14916), .c(n14911) );
no02f01  g9430 ( .o(n14918), .a(_net_10353), .b(n5710_1) );
no02f01  g9431 ( .o(n14919), .a(n9090), .b(n14918) );
oa12f01  g9432 ( .o(n14920), .a(n14919), .b(n9099), .c(n9088) );
no03f01  g9433 ( .o(n14921), .a(n14919), .b(n9099), .c(n9088) );
no02f01  g9434 ( .o(n14922), .a(n14921), .b(n8184) );
na02f01  g9435 ( .o(n14923), .a(n14922), .b(n14920) );
no02f01  g9436 ( .o(n14924), .a(n9132), .b(_net_10353) );
no02f01  g9437 ( .o(n14925), .a(n14924), .b(n9134) );
ao22f01  g9438 ( .o(n14926), .a(n14925), .b(n8200_1), .c(n8202), .d(_net_10353) );
na02f01  g9439 ( .o(n8697), .a(n14926), .b(n14923) );
no02f01  g9440 ( .o(n14928), .a(net_9157), .b(net_9156) );
no02f01  g9441 ( .o(n14929), .a(n10342), .b(n9168) );
no02f01  g9442 ( .o(n14930), .a(n14929), .b(n14928) );
na02f01  g9443 ( .o(n14931), .a(n14930), .b(n11392) );
in01f01  g9444 ( .o(n14932), .a(n14930) );
na02f01  g9445 ( .o(n14933), .a(n14932), .b(n11393) );
na03f01  g9446 ( .o(n14934), .a(n14933), .b(n14931), .c(n8638) );
ao12f01  g9447 ( .o(n14935), .a(n7883), .b(n8637), .c(_net_9315) );
na02f01  g9448 ( .o(n8702), .a(n14935), .b(n14934) );
in01f01  g9449 ( .o(n14937), .a(n14034) );
no02f01  g9450 ( .o(n14938), .a(n14937), .b(n9175) );
no02f01  g9451 ( .o(n14939), .a(n14034), .b(_net_10266) );
oa12f01  g9452 ( .o(n14940), .a(n6177_1), .b(n14939), .c(n14938) );
no02f01  g9453 ( .o(n14941), .a(n14039), .b(n9175) );
ao12f01  g9454 ( .o(n14942), .a(_net_10266), .b(n6945), .c(n9185) );
no03f01  g9455 ( .o(n14943), .a(n14942), .b(n14941), .c(n6846_1) );
ao12f01  g9456 ( .o(n14944), .a(n14943), .b(n6168), .c(_net_10266) );
na02f01  g9457 ( .o(n8707), .a(n14944), .b(n14940) );
ao22f01  g9458 ( .o(n14946), .a(n5842), .b(net_9756), .c(n5841), .d(net_192) );
na02f01  g9459 ( .o(n14947), .a(n5847), .b(net_10053) );
ao22f01  g9460 ( .o(n14948), .a(n5850), .b(net_9855), .c(n5849_1), .d(net_9954) );
na03f01  g9461 ( .o(n8712), .a(n14948), .b(n14947), .c(n14946) );
in01f01  g9462 ( .o(n14950), .a(_net_10108) );
ao12f01  g9463 ( .o(n14951), .a(n5658), .b(n6160_1), .c(x5289) );
oa12f01  g9464 ( .o(n8717), .a(n14951), .b(n6159), .c(n14950) );
na02f01  g9465 ( .o(n14953), .a(n8941), .b(_net_10331) );
na02f01  g9466 ( .o(n8722), .a(n14953), .b(n8943) );
ao12f01  g9467 ( .o(n14955), .a(n5658), .b(n7844), .c(_net_261) );
ao22f01  g9468 ( .o(n14956), .a(n7847), .b(x3949), .c(n7846), .d(net_9823) );
na02f01  g9469 ( .o(n8727), .a(n14956), .b(n14955) );
in01f01  g9470 ( .o(n14958), .a(_net_10308) );
ao12f01  g9471 ( .o(n14959), .a(n5658), .b(n5774), .c(x5901) );
oa12f01  g9472 ( .o(n8732), .a(n14959), .b(n5770), .c(n14958) );
na03f01  g9473 ( .o(n8737), .a(n13050), .b(n5884), .c(n5889) );
no02f01  g9474 ( .o(n14962), .a(n8126), .b(n13383) );
in01f01  g9475 ( .o(n14963), .a(n14962) );
no02f01  g9476 ( .o(n14964), .a(n14963), .b(n8131) );
na02f01  g9477 ( .o(n14965), .a(n14963), .b(n8131) );
na02f01  g9478 ( .o(n14966), .a(n14965), .b(n10948) );
no02f01  g9479 ( .o(n14967), .a(n8140_1), .b(_net_10154) );
no02f01  g9480 ( .o(n14968), .a(n8141), .b(n7778_1) );
no03f01  g9481 ( .o(n14969), .a(n14968), .b(n14967), .c(n10398) );
ao12f01  g9482 ( .o(n14970), .a(n14969), .b(n6760), .c(_net_10154) );
oa12f01  g9483 ( .o(n8742), .a(n14970), .b(n14966), .c(n14964) );
no02f01  g9484 ( .o(n14972), .a(_net_10365), .b(n7017_1) );
no02f01  g9485 ( .o(n14973), .a(n14972), .b(n7016) );
in01f01  g9486 ( .o(n14974), .a(n14973) );
na02f01  g9487 ( .o(n14975), .a(n7036), .b(n7020) );
na02f01  g9488 ( .o(n14976), .a(n14975), .b(n14974) );
na03f01  g9489 ( .o(n14977), .a(n14973), .b(n7036), .c(n7020) );
na02f01  g9490 ( .o(n8747), .a(n14977), .b(n14976) );
ao12f01  g9491 ( .o(n14979), .a(n5658), .b(n7844), .c(net_262) );
ao22f01  g9492 ( .o(n14980), .a(n7847), .b(x3889), .c(n7846), .d(net_9824) );
na02f01  g9493 ( .o(n8757), .a(n14980), .b(n14979) );
ao12f01  g9494 ( .o(n14982), .a(n5658), .b(n6160_1), .c(x4209) );
oa12f01  g9495 ( .o(n8767), .a(n14982), .b(n6159), .c(n7761) );
in01f01  g9496 ( .o(n14984), .a(_net_9644) );
no04f01  g9497 ( .o(n14985), .a(n8751), .b(n8749), .c(n7966), .d(n14984) );
no02f01  g9498 ( .o(n14986), .a(n8752), .b(n14984) );
oa12f01  g9499 ( .o(n14987), .a(_net_9641), .b(n14986), .c(n14816) );
na02f01  g9500 ( .o(n14988), .a(n9545), .b(_net_9644) );
oa22f01  g9501 ( .o(n14989), .a(n14988), .b(n8773), .c(n9791), .d(n14984) );
ao12f01  g9502 ( .o(n14990), .a(n14989), .b(n9495), .c(_net_9644) );
oa12f01  g9503 ( .o(n14991), .a(n14990), .b(n14987), .c(n9490) );
oa12f01  g9504 ( .o(n14992), .a(x6599), .b(n14991), .c(n14985) );
no02f01  g9505 ( .o(n8772), .a(n14992), .b(n2827) );
ao12f01  g9506 ( .o(n14994), .a(n7553), .b(n6028_1), .c(n6614_1) );
oa12f01  g9507 ( .o(n8777), .a(n14994), .b(n6022), .c(n7554) );
na02f01  g9508 ( .o(n14996), .a(n6056), .b(net_239) );
na02f01  g9509 ( .o(n14997), .a(n6055), .b(net_9967) );
ao22f01  g9510 ( .o(n14998), .a(n6062_1), .b(x5601), .c(n6060), .d(_net_10418) );
na04f01  g9511 ( .o(n8782), .a(n14998), .b(n14997), .c(n14996), .d(n6058) );
no02f01  g9512 ( .o(n15000), .a(n8173), .b(n8162) );
no02f01  g9513 ( .o(n15001), .a(_net_10365), .b(_net_9929) );
no02f01  g9514 ( .o(n15002), .a(n8164), .b(n15001) );
in01f01  g9515 ( .o(n15003), .a(n15002) );
ao12f01  g9516 ( .o(n15004), .a(n8184), .b(n15003), .c(n15000) );
oa12f01  g9517 ( .o(n15005), .a(n15004), .b(n15003), .c(n15000) );
oa12f01  g9518 ( .o(n15006), .a(_net_10365), .b(n8188), .c(_net_10364) );
ao12f01  g9519 ( .o(n15007), .a(n9144), .b(n15006), .c(n8190_1) );
ao12f01  g9520 ( .o(n15008), .a(n15007), .b(n8202), .c(_net_10365) );
na02f01  g9521 ( .o(n8787), .a(n15008), .b(n15005) );
no02f01  g9522 ( .o(n15010), .a(n5660), .b(n10694) );
ao22f01  g9523 ( .o(n15011), .a(n15010), .b(n6558), .c(n6577), .d(net_9689) );
ao22f01  g9524 ( .o(n15012), .a(n6606), .b(_net_9950), .c(n6599_1), .d(_net_9851) );
ao22f01  g9525 ( .o(n15013), .a(n6603), .b(net_10494), .c(n6572), .d(net_10389) );
na02f01  g9526 ( .o(n15014), .a(n6580), .b(net_9820) );
ao22f01  g9527 ( .o(n15015), .a(n6605), .b(net_10284), .c(n6585), .d(net_9721) );
na02f01  g9528 ( .o(n15016), .a(n15015), .b(n15014) );
na02f01  g9529 ( .o(n15017), .a(n6555), .b(net_9986) );
na02f01  g9530 ( .o(n15018), .a(n6573), .b(net_9887) );
na02f01  g9531 ( .o(n15019), .a(n6584_1), .b(net_9788) );
na02f01  g9532 ( .o(n15020), .a(n6592), .b(net_10179) );
na04f01  g9533 ( .o(n15021), .a(n15020), .b(n15019), .c(n15018), .d(n15017) );
na02f01  g9534 ( .o(n15022), .a(n6582), .b(net_9919) );
na02f01  g9535 ( .o(n15023), .a(n6602), .b(net_10018) );
ao22f01  g9536 ( .o(n15024), .a(n6597), .b(_net_9752), .c(n6590), .d(_net_10049) );
na03f01  g9537 ( .o(n15025), .a(n15024), .b(n15023), .c(n15022) );
no03f01  g9538 ( .o(n15026), .a(n15025), .b(n15021), .c(n15016) );
na04f01  g9539 ( .o(n8792), .a(n15026), .b(n15013), .c(n15012), .d(n15011) );
na02f01  g9540 ( .o(n15028), .a(n6038), .b(net_242) );
na02f01  g9541 ( .o(n15029), .a(n6037_1), .b(net_9871) );
ao22f01  g9542 ( .o(n15030), .a(n6044), .b(x5427), .c(n6042_1), .d(_net_10316) );
na04f01  g9543 ( .o(n8796), .a(n15030), .b(n15029), .c(n15028), .d(n6040) );
in01f01  g9544 ( .o(n15032), .a(_net_10534) );
oa22f01  g9545 ( .o(n8804), .a(n10629), .b(n15032), .c(n10685), .d(n5658) );
no02f01  g9546 ( .o(n15034), .a(n7804), .b(n7768_1) );
in01f01  g9547 ( .o(n15035), .a(n15034) );
na02f01  g9548 ( .o(n15036), .a(n15035), .b(n7791) );
na02f01  g9549 ( .o(n15037), .a(n15034), .b(n7792_1) );
na02f01  g9550 ( .o(n8809), .a(n15037), .b(n15036) );
na02f01  g9551 ( .o(n15039), .a(n7358), .b(_net_231) );
na02f01  g9552 ( .o(n15040), .a(n7352), .b(net_9662) );
ao22f01  g9553 ( .o(n15041), .a(n7357), .b(_net_10095), .c(n7353), .d(x6102) );
na04f01  g9554 ( .o(n8814), .a(n15041), .b(n15040), .c(n15039), .d(n7355_1) );
ao12f01  g9555 ( .o(n15043), .a(n5658), .b(n5678), .c(_net_254) );
ao22f01  g9556 ( .o(n15044), .a(n5681_1), .b(x4520), .c(n5680), .d(net_9717) );
na02f01  g9557 ( .o(n8819), .a(n15044), .b(n15043) );
na03f01  g9558 ( .o(n15046), .a(n5722), .b(n14279), .c(n5707) );
na04f01  g9559 ( .o(n15047), .a(n5705_1), .b(n5706), .c(n5721), .d(n8363_1) );
na04f01  g9560 ( .o(n15048), .a(n5711), .b(n5710_1), .c(n5719_1), .d(n5718) );
no03f01  g9561 ( .o(n15049), .a(n15048), .b(n15047), .c(n15046) );
ao12f01  g9562 ( .o(n8824), .a(n15049), .b(n10142), .c(n10140) );
oa22f01  g9563 ( .o(n8829), .a(n5694), .b(n5722), .c(n5692), .d(n5618) );
oa22f01  g9564 ( .o(n8834), .a(n5907), .b(n7871_1), .c(n5905), .d(n5537_1) );
oa22f01  g9565 ( .o(n8839), .a(n7367), .b(n10379), .c(n7365_1), .d(n5649) );
no02f01  g9566 ( .o(n15054), .a(n10977), .b(n12072) );
oa12f01  g9567 ( .o(n15055), .a(n10948), .b(n10978), .c(_net_10150) );
na02f01  g9568 ( .o(n15056), .a(n10992), .b(n12072) );
no02f01  g9569 ( .o(n15057), .a(n11160), .b(n10398) );
ao22f01  g9570 ( .o(n15058), .a(n15057), .b(n15056), .c(n6760), .d(_net_10150) );
oa12f01  g9571 ( .o(n8844), .a(n15058), .b(n15055), .c(n15054) );
in01f01  g9572 ( .o(n15060), .a(_net_10317) );
ao12f01  g9573 ( .o(n15061), .a(n5658), .b(n5774), .c(x5364) );
oa12f01  g9574 ( .o(n8857), .a(n15061), .b(n5770), .c(n15060) );
ao12f01  g9575 ( .o(n15063), .a(n5658), .b(n6887), .c(x4520) );
oa12f01  g9576 ( .o(n8862), .a(n15063), .b(n6885_1), .c(n9200) );
no02f01  g9577 ( .o(n15065), .a(n9111), .b(n9083) );
in01f01  g9578 ( .o(n15066), .a(n15065) );
ao12f01  g9579 ( .o(n15067), .a(n15066), .b(n9108), .c(n9102) );
na02f01  g9580 ( .o(n15068), .a(n9108), .b(n9102) );
oa12f01  g9581 ( .o(n15069), .a(n8183), .b(n15065), .c(n15068) );
na02f01  g9582 ( .o(n15070), .a(n9137), .b(n9110) );
no02f01  g9583 ( .o(n15071), .a(n9138), .b(n9144) );
ao22f01  g9584 ( .o(n15072), .a(n15071), .b(n15070), .c(n8202), .d(_net_10356) );
oa12f01  g9585 ( .o(n8867), .a(n15072), .b(n15069), .c(n15067) );
na02f01  g9586 ( .o(n15074), .a(_net_10324), .b(n7029) );
na02f01  g9587 ( .o(n8872), .a(n15074), .b(n9781) );
bf01f01  g9588 ( .o(x19), .a(x185142) );
bf01f01  g9589 ( .o(x916), .a(x185142) );
bf01f01  g9590 ( .o(x936), .a(x185142) );
bf01f01  g9591 ( .o(x948), .a(x185142) );
bf01f01  g9592 ( .o(x921), .a(x185142) );
bf01f01  g9593 ( .o(x957), .a(x185142) );
bf01f01  g9594 ( .o(x906), .a(x185142) );
bf01f01  g9595 ( .o(x472), .a(_net_8847) );
bf01f01  g9596 ( .o(x941), .a(x185142) );
bf01f01  g9597 ( .o(x926), .a(x185142) );
bf01f01  g9598 ( .o(x813), .a(x6599) );
bf01f01  g9599 ( .o(x911), .a(x185142) );
bf01f01  g9600 ( .o(x898), .a(x185142) );
bf01f01  g9601 ( .o(x890), .a(x185142) );
bf01f01  g9602 ( .o(x931), .a(x185142) );
bf01f01  g9603 ( .o(n510), .a(net_9141) );
bf01f01  g9604 ( .o(n524), .a(net_9337) );
bf01f01  g9605 ( .o(n558), .a(net_10408) );
bf01f01  g9606 ( .o(n628), .a(net_92) );
bf01f01  g9607 ( .o(n638), .a(net_9461) );
bf01f01  g9608 ( .o(n657), .a(net_9328) );
bf01f01  g9609 ( .o(n721), .a(net_9281) );
bf01f01  g9610 ( .o(n736), .a(net_9260) );
bf01f01  g9611 ( .o(n746), .a(net_9163) );
bf01f01  g9612 ( .o(n751), .a(net_287) );
bf01f01  g9613 ( .o(n770), .a(net_9463) );
bf01f01  g9614 ( .o(n774), .a(net_284) );
bf01f01  g9615 ( .o(n917), .a(x2165) );
bf01f01  g9616 ( .o(n932), .a(net_9466) );
bf01f01  g9617 ( .o(n940), .a(x3606) );
bf01f01  g9618 ( .o(n945), .a(net_9284) );
bf01f01  g9619 ( .o(n958), .a(x2400) );
bf01f01  g9620 ( .o(n968), .a(_net_9502) );
bf01f01  g9621 ( .o(n978), .a(net_307) );
bf01f01  g9622 ( .o(n987), .a(_net_9160) );
bf01f01  g9623 ( .o(n992), .a(net_108) );
bf01f01  g9624 ( .o(n1107), .a(net_281) );
bf01f01  g9625 ( .o(n1121), .a(net_310) );
bf01f01  g9626 ( .o(n1175), .a(net_10518) );
bf01f01  g9627 ( .o(n1218), .a(net_9132) );
bf01f01  g9628 ( .o(n1237), .a(net_10303) );
bf01f01  g9629 ( .o(n1282), .a(_net_10244) );
bf01f01  g9630 ( .o(n1296), .a(_net_9258) );
bf01f01  g9631 ( .o(n1310), .a(x2098) );
bf01f01  g9632 ( .o(n1335), .a(net_9454) );
bf01f01  g9633 ( .o(n1364), .a(net_9584) );
bf01f01  g9634 ( .o(n1388), .a(net_9281) );
bf01f01  g9635 ( .o(n1397), .a(net_9286) );
bf01f01  g9636 ( .o(n1411), .a(net_9147) );
bf01f01  g9637 ( .o(n1440), .a(net_299) );
bf01f01  g9638 ( .o(n1474), .a(net_9148) );
bf01f01  g9639 ( .o(n1488), .a(net_9338) );
bf01f01  g9640 ( .o(n1517), .a(net_305) );
bf01f01  g9641 ( .o(n1536), .a(net_9330) );
bf01f01  g9642 ( .o(n1545), .a(net_9456) );
bf01f01  g9643 ( .o(n1579), .a(net_9137) );
bf01f01  g9644 ( .o(n1582), .a(x3314) );
bf01f01  g9645 ( .o(n1602), .a(net_311) );
bf01f01  g9646 ( .o(n1605), .a(net_9127) );
bf01f01  g9647 ( .o(n1618), .a(net_116) );
bf01f01  g9648 ( .o(n1623), .a(net_9303) );
bf01f01  g9649 ( .o(n1627), .a(net_302) );
bf01f01  g9650 ( .o(n1661), .a(net_9288) );
bf01f01  g9651 ( .o(n1715), .a(x1459) );
bf01f01  g9652 ( .o(n1735), .a(net_9451) );
bf01f01  g9653 ( .o(n1783), .a(x3360) );
bf01f01  g9654 ( .o(n1826), .a(x2707) );
bf01f01  g9655 ( .o(n1831), .a(net_9136) );
bf01f01  g9656 ( .o(n1839), .a(x3558) );
bf01f01  g9657 ( .o(n1863), .a(x3071) );
bf01f01  g9658 ( .o(n1872), .a(x2589) );
bf01f01  g9659 ( .o(n1881), .a(net_9182) );
bf01f01  g9660 ( .o(n2070), .a(net_9116) );
bf01f01  g9661 ( .o(n2130), .a(_net_10434) );
bf01f01  g9662 ( .o(n2140), .a(net_9151) );
bf01f01  g9663 ( .o(n2160), .a(_net_10543) );
bf01f01  g9664 ( .o(n2169), .a(x3565) );
bf01f01  g9665 ( .o(n2189), .a(net_9146) );
bf01f01  g9666 ( .o(n2202), .a(net_10408) );
bf01f01  g9667 ( .o(n2217), .a(net_9582) );
bf01f01  g9668 ( .o(n2246), .a(_net_10543) );
bf01f01  g9669 ( .o(n2325), .a(x3534) );
bf01f01  g9670 ( .o(n2334), .a(net_9134) );
bf01f01  g9671 ( .o(n2338), .a(net_282) );
bf01f01  g9672 ( .o(n2367), .a(net_136) );
bf01f01  g9673 ( .o(n2371), .a(x555) );
bf01f01  g9674 ( .o(n2404), .a(net_9158) );
bf01f01  g9675 ( .o(n2414), .a(net_9659) );
bf01f01  g9676 ( .o(n2449), .a(net_139) );
bf01f01  g9677 ( .o(n2453), .a(x2214) );
bf01f01  g9678 ( .o(n2473), .a(net_9305) );
bf01f01  g9679 ( .o(n2497), .a(net_9184) );
bf01f01  g9680 ( .o(n2532), .a(net_98) );
bf01f01  g9681 ( .o(n2537), .a(net_9452) );
bf01f01  g9682 ( .o(n2560), .a(x480) );
bf01f01  g9683 ( .o(n2568), .a(x798) );
bf01f01  g9684 ( .o(n2647), .a(_net_10535) );
bf01f01  g9685 ( .o(n2662), .a(_net_9267) );
bf01f01  g9686 ( .o(n2685), .a(net_9154) );
bf01f01  g9687 ( .o(n2720), .a(_net_9646) );
bf01f01  g9688 ( .o(n2769), .a(x1865) );
bf01f01  g9689 ( .o(n2798), .a(x2477) );
bf01f01  g9690 ( .o(n2817), .a(x1743) );
bf01f01  g9691 ( .o(n2832), .a(net_9438) );
bf01f01  g9692 ( .o(n2851), .a(net_9333) );
bf01f01  g9693 ( .o(n2908), .a(net_9439) );
bf01f01  g9694 ( .o(n2942), .a(net_9441) );
bf01f01  g9695 ( .o(n2956), .a(net_10519) );
bf01f01  g9696 ( .o(n3034), .a(x1660) );
bf01f01  g9697 ( .o(n3039), .a(net_10516) );
bf01f01  g9698 ( .o(n3073), .a(net_285) );
bf01f01  g9699 ( .o(n3097), .a(net_296) );
bf01f01  g9700 ( .o(n3161), .a(net_138) );
bf01f01  g9701 ( .o(n3210), .a(net_114) );
bf01f01  g9702 ( .o(n3220), .a(_net_9118) );
bf01f01  g9703 ( .o(n3234), .a(net_9122) );
bf01f01  g9704 ( .o(n3247), .a(x1911) );
bf01f01  g9705 ( .o(n3291), .a(x3599) );
bf01f01  g9706 ( .o(n3310), .a(net_9157) );
bf01f01  g9707 ( .o(n3359), .a(net_9576) );
bf01f01  g9708 ( .o(n3413), .a(net_9459) );
bf01f01  g9709 ( .o(n3416), .a(net_9575) );
bf01f01  g9710 ( .o(n3426), .a(net_9446) );
bf01f01  g9711 ( .o(n3440), .a(net_10513) );
bf01f01  g9712 ( .o(n3495), .a(net_9140) );
bf01f01  g9713 ( .o(n3509), .a(net_9150) );
bf01f01  g9714 ( .o(n3623), .a(net_9259) );
bf01f01  g9715 ( .o(n3633), .a(_net_9266) );
bf01f01  g9716 ( .o(n3647), .a(x6599) );
bf01f01  g9717 ( .o(n3746), .a(net_10519) );
bf01f01  g9718 ( .o(n3754), .a(x3194) );
bf01f01  g9719 ( .o(n3758), .a(x3534) );
bf01f01  g9720 ( .o(n3782), .a(x3300) );
bf01f01  g9721 ( .o(n3792), .a(net_9468) );
bf01f01  g9722 ( .o(n3835), .a(net_309) );
bf01f01  g9723 ( .o(n3919), .a(net_9280) );
bf01f01  g9724 ( .o(n3933), .a(net_289) );
bf01f01  g9725 ( .o(n3937), .a(net_9152) );
bf01f01  g9726 ( .o(n3957), .a(net_147) );
bf01f01  g9727 ( .o(n3976), .a(x784) );
bf01f01  g9728 ( .o(n4084), .a(net_9283) );
bf01f01  g9729 ( .o(n4088), .a(net_9263) );
bf01f01  g9730 ( .o(n4108), .a(net_9453) );
bf01f01  g9731 ( .o(n4116), .a(net_9135) );
bf01f01  g9732 ( .o(n4120), .a(net_9340) );
bf01f01  g9733 ( .o(n4133), .a(net_10518) );
bf01f01  g9734 ( .o(n4151), .a(net_135) );
bf01f01  g9735 ( .o(n4215), .a(net_10198) );
bf01f01  g9736 ( .o(n4255), .a(net_301) );
bf01f01  g9737 ( .o(n4279), .a(_net_10349) );
bf01f01  g9738 ( .o(n4312), .a(net_9155) );
bf01f01  g9739 ( .o(n4316), .a(net_9578) );
bf01f01  g9740 ( .o(n4351), .a(net_143) );
bf01f01  g9741 ( .o(n4364), .a(net_9465) );
bf01f01  g9742 ( .o(n4368), .a(net_9126) );
bf01f01  g9743 ( .o(n4401), .a(_net_10543) );
bf01f01  g9744 ( .o(n4430), .a(net_9123) );
bf01f01  g9745 ( .o(n4463), .a(net_10513) );
bf01f01  g9746 ( .o(n4477), .a(x1598) );
bf01f01  g9747 ( .o(n4491), .a(x3507) );
bf01f01  g9748 ( .o(n4516), .a(_net_10329) );
bf01f01  g9749 ( .o(n4535), .a(net_306) );
bf01f01  g9750 ( .o(n4584), .a(net_95) );
bf01f01  g9751 ( .o(n4598), .a(net_9570) );
bf01f01  g9752 ( .o(n4627), .a(net_145) );
bf01f01  g9753 ( .o(n4647), .a(net_292) );
bf01f01  g9754 ( .o(n4650), .a(net_9128) );
bf01f01  g9755 ( .o(n4668), .a(net_9253) );
bf01f01  g9756 ( .o(n4682), .a(net_10198) );
bf01f01  g9757 ( .o(n4692), .a(net_295) );
bf01f01  g9758 ( .o(n4700), .a(net_9265) );
bf01f01  g9759 ( .o(n4724), .a(_net_10528) );
bf01f01  g9760 ( .o(n4784), .a(net_297) );
bf01f01  g9761 ( .o(n4793), .a(net_10541) );
bf01f01  g9762 ( .o(n4842), .a(net_9131) );
bf01f01  g9763 ( .o(n4861), .a(net_105) );
bf01f01  g9764 ( .o(n4875), .a(x3327) );
bf01f01  g9765 ( .o(n4904), .a(net_10517) );
bf01f01  g9766 ( .o(n4927), .a(x3653) );
bf01f01  g9767 ( .o(n4946), .a(net_10542) );
bf01f01  g9768 ( .o(n4976), .a(net_308) );
bf01f01  g9769 ( .o(n5038), .a(net_99) );
bf01f01  g9770 ( .o(n5052), .a(net_9234) );
bf01f01  g9771 ( .o(n5087), .a(net_9304) );
bf01f01  g9772 ( .o(n5101), .a(net_9282) );
bf01f01  g9773 ( .o(n5139), .a(net_9133) );
bf01f01  g9774 ( .o(n5147), .a(net_141) );
bf01f01  g9775 ( .o(n5157), .a(net_9445) );
bf01f01  g9776 ( .o(n5161), .a(net_9327) );
bf01f01  g9777 ( .o(n5165), .a(net_9464) );
bf01f01  g9778 ( .o(n5194), .a(net_304) );
bf01f01  g9779 ( .o(n5212), .a(x1547) );
bf01f01  g9780 ( .o(n5262), .a(net_298) );
bf01f01  g9781 ( .o(n5266), .a(net_9125) );
bf01f01  g9782 ( .o(n5279), .a(net_9139) );
bf01f01  g9783 ( .o(n5297), .a(x3320) );
bf01f01  g9784 ( .o(n5306), .a(x6599) );
bf01f01  g9785 ( .o(n5351), .a(net_9144) );
bf01f01  g9786 ( .o(n5370), .a(net_9156) );
bf01f01  g9787 ( .o(n5375), .a(net_9339) );
bf01f01  g9788 ( .o(n5403), .a(net_10536) );
bf01f01  g9789 ( .o(n5408), .a(net_9285) );
bf01f01  g9790 ( .o(n5431), .a(net_9255) );
bf01f01  g9791 ( .o(n5445), .a(net_9387) );
no03f01  g9792 ( .o(n5449), .a(n6461), .b(n5633), .c(n6354) );
bf01f01  g9793 ( .o(n5473), .a(net_9448) );
bf01f01  g9794 ( .o(n5477), .a(net_9329) );
bf01f01  g9795 ( .o(n5495), .a(net_9264) );
bf01f01  g9796 ( .o(n5504), .a(x3338) );
bf01f01  g9797 ( .o(n5508), .a(net_9284) );
bf01f01  g9798 ( .o(n5582), .a(net_288) );
bf01f01  g9799 ( .o(n5585), .a(x3613) );
bf01f01  g9800 ( .o(n5589), .a(x2333) );
bf01f01  g9801 ( .o(n5594), .a(net_290) );
bf01f01  g9802 ( .o(n5597), .a(x3307) );
bf01f01  g9803 ( .o(n5601), .a(net_9449) );
bf01f01  g9804 ( .o(n5614), .a(x1503) );
bf01f01  g9805 ( .o(n5629), .a(net_9469) );
bf01f01  g9806 ( .o(n5638), .a(net_9335) );
bf01f01  g9807 ( .o(n5651), .a(net_140) );
bf01f01  g9808 ( .o(n5681), .a(net_294) );
bf01f01  g9809 ( .o(n5714), .a(x2648) );
bf01f01  g9810 ( .o(n5777), .a(net_109) );
bf01f01  g9811 ( .o(n5812), .a(net_9336) );
bf01f01  g9812 ( .o(n5815), .a(_net_9502) );
bf01f01  g9813 ( .o(n5853), .a(net_9543) );
bf01f01  g9814 ( .o(n5917), .a(x3621) );
bf01f01  g9815 ( .o(n5935), .a(net_9283) );
bf01f01  g9816 ( .o(n5939), .a(net_9282) );
bf01f01  g9817 ( .o(n5974), .a(net_9138) );
bf01f01  g9818 ( .o(n5998), .a(net_9334) );
bf01f01  g9819 ( .o(n6001), .a(net_10516) );
bf01f01  g9820 ( .o(n6009), .a(net_9119) );
bf01f01  g9821 ( .o(n6067), .a(net_134) );
bf01f01  g9822 ( .o(n6091), .a(net_300) );
bf01f01  g9823 ( .o(n6095), .a(net_9462) );
bf01f01  g9824 ( .o(n6099), .a(net_9467) );
bf01f01  g9825 ( .o(n6102), .a(net_9252) );
bf01f01  g9826 ( .o(n6145), .a(net_107) );
bf01f01  g9827 ( .o(n6169), .a(net_9287) );
bf01f01  g9828 ( .o(n6177), .a(net_97) );
bf01f01  g9829 ( .o(n6181), .a(net_144) );
bf01f01  g9830 ( .o(n6235), .a(net_96) );
bf01f01  g9831 ( .o(n6240), .a(net_283) );
bf01f01  g9832 ( .o(n6254), .a(net_9129) );
bf01f01  g9833 ( .o(n6272), .a(x3349) );
bf01f01  g9834 ( .o(n6302), .a(net_9442) );
bf01f01  g9835 ( .o(n6360), .a(net_9331) );
bf01f01  g9836 ( .o(n6369), .a(net_9306) );
bf01f01  g9837 ( .o(n6401), .a(net_9262) );
bf01f01  g9838 ( .o(n6460), .a(x3249) );
bf01f01  g9839 ( .o(n6464), .a(x2826) );
bf01f01  g9840 ( .o(n6493), .a(x2027) );
bf01f01  g9841 ( .o(n6507), .a(x2767) );
bf01f01  g9842 ( .o(n6579), .a(x1974) );
bf01f01  g9843 ( .o(n6713), .a(x2968) );
bf01f01  g9844 ( .o(n6782), .a(net_9143) );
no02f01  g9845 ( .o(n6865), .a(n11966), .b(n6686) );
bf01f01  g9846 ( .o(n6910), .a(net_9120) );
bf01f01  g9847 ( .o(n6944), .a(net_115) );
bf01f01  g9848 ( .o(n6958), .a(net_9577) );
bf01f01  g9849 ( .o(n6962), .a(net_9583) );
bf01f01  g9850 ( .o(n6966), .a(x3133) );
bf01f01  g9851 ( .o(n6985), .a(net_9440) );
bf01f01  g9852 ( .o(n6993), .a(net_137) );
bf01f01  g9853 ( .o(n7007), .a(x3507) );
bf01f01  g9854 ( .o(n7021), .a(x6599) );
bf01f01  g9855 ( .o(n7030), .a(x3588) );
bf01f01  g9856 ( .o(n7044), .a(net_9455) );
bf01f01  g9857 ( .o(n7078), .a(net_291) );
bf01f01  g9858 ( .o(n7086), .a(net_9574) );
bf01f01  g9859 ( .o(n7095), .a(net_9257) );
bf01f01  g9860 ( .o(n7100), .a(net_9458) );
bf01f01  g9861 ( .o(n7108), .a(net_10093) );
bf01f01  g9862 ( .o(n7206), .a(net_10303) );
bf01f01  g9863 ( .o(n7270), .a(_net_10224) );
bf01f01  g9864 ( .o(n7304), .a(net_9130) );
bf01f01  g9865 ( .o(n7308), .a(_net_10139) );
bf01f01  g9866 ( .o(n7317), .a(net_9307) );
bf01f01  g9867 ( .o(n7355), .a(net_9153) );
bf01f01  g9868 ( .o(n7398), .a(net_9261) );
bf01f01  g9869 ( .o(n7436), .a(x1418) );
bf01f01  g9870 ( .o(n7480), .a(net_9450) );
bf01f01  g9871 ( .o(n7538), .a(x1792) );
bf01f01  g9872 ( .o(n7575), .a(x2531) );
bf01f01  g9873 ( .o(n7580), .a(net_112) );
bf01f01  g9874 ( .o(n7613), .a(net_9149) );
bf01f01  g9875 ( .o(n7617), .a(net_9444) );
bf01f01  g9876 ( .o(n7640), .a(x2890) );
bf01f01  g9877 ( .o(n7704), .a(net_106) );
bf01f01  g9878 ( .o(n7734), .a(net_286) );
bf01f01  g9879 ( .o(n7782), .a(net_9254) );
bf01f01  g9880 ( .o(n7830), .a(net_9124) );
bf01f01  g9881 ( .o(n7862), .a(net_303) );
bf01f01  g9882 ( .o(n7885), .a(net_142) );
bf01f01  g9883 ( .o(n7902), .a(net_9159) );
no04f01  g9884 ( .o(n7906), .a(n13308), .b(n13307), .c(n13306), .d(n7976) );
bf01f01  g9885 ( .o(n7925), .a(net_94) );
bf01f01  g9886 ( .o(n7954), .a(net_9457) );
bf01f01  g9887 ( .o(n7957), .a(net_9285) );
bf01f01  g9888 ( .o(n7992), .a(_net_9244) );
bf01f01  g9889 ( .o(n8055), .a(net_146) );
bf01f01  g9890 ( .o(n8063), .a(net_9579) );
bf01f01  g9891 ( .o(n8067), .a(x3022) );
bf01f01  g9892 ( .o(n8076), .a(net_93) );
bf01f01  g9893 ( .o(n8120), .a(net_9287) );
bf01f01  g9894 ( .o(n8210), .a(_net_10454) );
bf01f01  g9895 ( .o(n8219), .a(net_9447) );
bf01f01  g9896 ( .o(n8227), .a(net_9121) );
bf01f01  g9897 ( .o(n8235), .a(net_9256) );
bf01f01  g9898 ( .o(n8264), .a(net_10517) );
bf01f01  g9899 ( .o(n8272), .a(net_9142) );
bf01f01  g9900 ( .o(n8305), .a(x6599) );
bf01f01  g9901 ( .o(n8339), .a(_net_9646) );
bf01f01  g9902 ( .o(n8368), .a(net_293) );
bf01f01  g9903 ( .o(n8376), .a(net_9286) );
bf01f01  g9904 ( .o(n8380), .a(x3574) );
bf01f01  g9905 ( .o(n8433), .a(net_9280) );
bf01f01  g9906 ( .o(n8443), .a(net_9342) );
bf01f01  g9907 ( .o(n8486), .a(x2278) );
bf01f01  g9908 ( .o(n8501), .a(net_9443) );
bf01f01  g9909 ( .o(n8529), .a(_net_9378) );
bf01f01  g9910 ( .o(n8562), .a(net_9251) );
bf01f01  g9911 ( .o(n8577), .a(_net_9606) );
bf01f01  g9912 ( .o(n8646), .a(net_312) );
bf01f01  g9913 ( .o(n8693), .a(net_9332) );
bf01f01  g9914 ( .o(n8800), .a(x732) );
bf01f01  g9915 ( .o(n8849), .a(net_9460) );
bf01f01  g9916 ( .o(n8853), .a(net_9341) );
bf01f01  g9917 ( .o(n8876), .a(net_9145) );
ms00f80  l0001 ( .o(net_9715), .ck(clk), .d(n500) );
ms00f80  l0002 ( .o(net_9939), .ck(clk), .d(n505) );
ms00f80  l0003 ( .o(x1170), .ck(clk), .d(n510) );
ms00f80  l0004 ( .o(_net_9400), .ck(clk), .d(n514) );
ms00f80  l0005 ( .o(net_9956), .ck(clk), .d(n519) );
ms00f80  l0006 ( .o(net_9337), .ck(clk), .d(n524) );
ms00f80  l0007 ( .o(_net_9414), .ck(clk), .d(n528) );
ms00f80  l0008 ( .o(_net_10136), .ck(clk), .d(n533) );
ms00f80  l0009 ( .o(_net_10312), .ck(clk), .d(n538) );
ms00f80  l0010 ( .o(net_116), .ck(clk), .d(n543) );
ms00f80  l0011 ( .o(net_9538), .ck(clk), .d(n548) );
ms00f80  l0012 ( .o(net_9940), .ck(clk), .d(n553) );
ms00f80  l0013 ( .o(_net_10348), .ck(clk), .d(n558) );
ms00f80  l0014 ( .o(_net_10029), .ck(clk), .d(n563) );
ms00f80  l0015 ( .o(net_10299), .ck(clk), .d(n568) );
ms00f80  l0016 ( .o(net_197), .ck(clk), .d(n573) );
ms00f80  l0017 ( .o(_net_9589), .ck(clk), .d(n578) );
ms00f80  l0018 ( .o(net_9869), .ck(clk), .d(n583) );
ms00f80  l0019 ( .o(net_9990), .ck(clk), .d(n588) );
ms00f80  l0020 ( .o(_net_9371), .ck(clk), .d(n593) );
ms00f80  l0021 ( .o(net_10065), .ck(clk), .d(n598) );
ms00f80  l0022 ( .o(_net_10104), .ck(clk), .d(n603) );
ms00f80  l0023 ( .o(_net_10258), .ck(clk), .d(n608) );
ms00f80  l0024 ( .o(_net_278), .ck(clk), .d(n613) );
ms00f80  l0025 ( .o(_net_9272), .ck(clk), .d(n618) );
ms00f80  l0026 ( .o(_net_9238), .ck(clk), .d(n623) );
ms00f80  l0027 ( .o(net_10520), .ck(clk), .d(n628) );
ms00f80  l0028 ( .o(net_10007), .ck(clk), .d(n633) );
ms00f80  l0029 ( .o(net_9461), .ck(clk), .d(n638) );
ms00f80  l0030 ( .o(net_9619), .ck(clk), .d(n642) );
ms00f80  l0031 ( .o(net_9135), .ck(clk), .d(n647) );
ms00f80  l0032 ( .o(net_9583), .ck(clk), .d(n652) );
ms00f80  l0033 ( .o(net_9328), .ck(clk), .d(n657) );
ms00f80  l0034 ( .o(_net_10137), .ck(clk), .d(n661) );
ms00f80  l0035 ( .o(net_9206), .ck(clk), .d(n666) );
ms00f80  l0036 ( .o(_net_10110), .ck(clk), .d(n671) );
ms00f80  l0037 ( .o(_net_10429), .ck(clk), .d(n676) );
ms00f80  l0038 ( .o(_net_10144), .ck(clk), .d(n681) );
ms00f80  l0039 ( .o(_net_8825), .ck(clk), .d(n686) );
ms00f80  l0040 ( .o(_net_10256), .ck(clk), .d(n691) );
ms00f80  l0041 ( .o(_net_9249), .ck(clk), .d(n696) );
ms00f80  l0042 ( .o(net_9921), .ck(clk), .d(n701) );
ms00f80  l0043 ( .o(_net_10219), .ck(clk), .d(n706) );
ms00f80  l0044 ( .o(net_10034), .ck(clk), .d(n711) );
ms00f80  l0045 ( .o(net_9867), .ck(clk), .d(n716) );
ms00f80  l0046 ( .o(net_9505), .ck(clk), .d(n721) );
ms00f80  l0047 ( .o(net_9917), .ck(clk), .d(n726) );
ms00f80  l0048 ( .o(_net_10323), .ck(clk), .d(n731) );
ms00f80  l0049 ( .o(_net_9554), .ck(clk), .d(n736) );
ms00f80  l0050 ( .o(_net_10264), .ck(clk), .d(n741) );
ms00f80  l0051 ( .o(_net_9164), .ck(clk), .d(n746) );
ms00f80  l0052 ( .o(net_287), .ck(clk), .d(n751) );
ms00f80  l0053 ( .o(net_9130), .ck(clk), .d(n755) );
ms00f80  l0054 ( .o(net_9748), .ck(clk), .d(n760) );
ms00f80  l0055 ( .o(_net_10139), .ck(clk), .d(n765) );
ms00f80  l0056 ( .o(net_9463), .ck(clk), .d(n770) );
ms00f80  l0057 ( .o(net_284), .ck(clk), .d(n774) );
ms00f80  l0058 ( .o(_net_8831), .ck(clk), .d(n778) );
ms00f80  l0059 ( .o(net_10088), .ck(clk), .d(n783) );
ms00f80  l0060 ( .o(_net_10216), .ck(clk), .d(n788) );
ms00f80  l0061 ( .o(net_8822), .ck(clk), .d(n793) );
ms00f80  l0062 ( .o(_net_9591), .ck(clk), .d(n798) );
ms00f80  l0063 ( .o(_net_10205), .ck(clk), .d(n803) );
ms00f80  l0064 ( .o(net_9986), .ck(clk), .d(n808) );
ms00f80  l0065 ( .o(net_9897), .ck(clk), .d(n813) );
ms00f80  l0066 ( .o(_net_9362), .ck(clk), .d(n818) );
ms00f80  l0067 ( .o(net_9669), .ck(clk), .d(n823) );
ms00f80  l0068 ( .o(_net_10431), .ck(clk), .d(n828) );
ms00f80  l0069 ( .o(net_9749), .ck(clk), .d(n833) );
ms00f80  l0070 ( .o(_net_10478), .ck(clk), .d(n838) );
ms00f80  l0071 ( .o(net_9724), .ck(clk), .d(n843) );
ms00f80  l0072 ( .o(_net_185), .ck(clk), .d(n848) );
ms00f80  l0073 ( .o(net_10502), .ck(clk), .d(n853) );
ms00f80  l0074 ( .o(_net_131), .ck(clk), .d(n858) );
ms00f80  l0075 ( .o(net_9687), .ck(clk), .d(n863) );
ms00f80  l0076 ( .o(_net_9831), .ck(clk), .d(n868) );
ms00f80  l0077 ( .o(_net_9247), .ck(clk), .d(n873) );
ms00f80  l0078 ( .o(net_246), .ck(clk), .d(n878) );
ms00f80  l0079 ( .o(net_9133), .ck(clk), .d(n883) );
ms00f80  l0080 ( .o(_net_9202), .ck(clk), .d(n888) );
ms00f80  l0081 ( .o(net_9208), .ck(clk), .d(n893) );
ms00f80  l0082 ( .o(net_10005), .ck(clk), .d(n898) );
ms00f80  l0083 ( .o(net_9616), .ck(clk), .d(n903) );
ms00f80  l0084 ( .o(net_10450), .ck(clk), .d(n908) );
ms00f80  l0085 ( .o(_net_10248), .ck(clk), .d(n913) );
ms00f80  l0086 ( .o(net_9488), .ck(clk), .d(n917) );
ms00f80  l0087 ( .o(_net_10203), .ck(clk), .d(n922) );
ms00f80  l0088 ( .o(_net_122), .ck(clk), .d(n927) );
ms00f80  l0089 ( .o(net_9466), .ck(clk), .d(n932) );
ms00f80  l0090 ( .o(net_9229), .ck(clk), .d(n936) );
ms00f80  l0091 ( .o(net_9154), .ck(clk), .d(n940) );
ms00f80  l0092 ( .o(net_9284), .ck(clk), .d(n945) );
ms00f80  l0093 ( .o(_net_269), .ck(clk), .d(n949) );
ms00f80  l0094 ( .o(_net_9834), .ck(clk), .d(n954) );
ms00f80  l0095 ( .o(net_9484), .ck(clk), .d(n958) );
ms00f80  l0096 ( .o(net_9880), .ck(clk), .d(n963) );
ms00f80  l0097 ( .o(net_9543), .ck(clk), .d(n968) );
ms00f80  l0098 ( .o(net_9618), .ck(clk), .d(n973) );
ms00f80  l0099 ( .o(net_307), .ck(clk), .d(n978) );
ms00f80  l0100 ( .o(_net_9160), .ck(clk), .d(n982) );
ms00f80  l0101 ( .o(_net_10092), .ck(clk), .d(n987) );
ms00f80  l0102 ( .o(net_239), .ck(clk), .d(n992) );
ms00f80  l0103 ( .o(net_9604), .ck(clk), .d(n997) );
ms00f80  l0104 ( .o(_net_9346), .ck(clk), .d(n1002) );
ms00f80  l0105 ( .o(net_9175), .ck(clk), .d(n1007) );
ms00f80  l0106 ( .o(net_217), .ck(clk), .d(n1012) );
ms00f80  l0107 ( .o(net_9994), .ck(clk), .d(n1017) );
ms00f80  l0108 ( .o(net_8838), .ck(clk), .d(n1022) );
ms00f80  l0109 ( .o(_net_9581), .ck(clk), .d(n1027) );
ms00f80  l0110 ( .o(_net_8839), .ck(clk), .d(n1032) );
ms00f80  l0111 ( .o(_net_119), .ck(clk), .d(n1037) );
ms00f80  l0112 ( .o(net_9818), .ck(clk), .d(n1042) );
ms00f80  l0113 ( .o(_net_9237), .ck(clk), .d(n1047) );
ms00f80  l0114 ( .o(net_9712), .ck(clk), .d(n1052) );
ms00f80  l0115 ( .o(_net_10470), .ck(clk), .d(n1057) );
ms00f80  l0116 ( .o(_net_9325), .ck(clk), .d(n1062) );
ms00f80  l0117 ( .o(net_9694), .ck(clk), .d(n1067) );
ms00f80  l0118 ( .o(net_9774), .ck(clk), .d(n1072) );
ms00f80  l0119 ( .o(net_9678), .ck(clk), .d(n1077) );
ms00f80  l0120 ( .o(net_141), .ck(clk), .d(n1082) );
ms00f80  l0121 ( .o(net_10179), .ck(clk), .d(n1087) );
ms00f80  l0122 ( .o(_net_9518), .ck(clk), .d(n1092) );
ms00f80  l0123 ( .o(net_135), .ck(clk), .d(n1097) );
ms00f80  l0124 ( .o(_net_10116), .ck(clk), .d(n1102) );
ms00f80  l0125 ( .o(net_281), .ck(clk), .d(n1107) );
ms00f80  l0126 ( .o(net_9790), .ck(clk), .d(n1111) );
ms00f80  l0127 ( .o(_net_9188), .ck(clk), .d(n1116) );
ms00f80  l0128 ( .o(net_310), .ck(clk), .d(n1121) );
ms00f80  l0129 ( .o(_net_9192), .ck(clk), .d(n1125) );
ms00f80  l0130 ( .o(_net_9729), .ck(clk), .d(n1130) );
ms00f80  l0131 ( .o(net_9821), .ck(clk), .d(n1135) );
ms00f80  l0132 ( .o(net_9122), .ck(clk), .d(n1140) );
ms00f80  l0133 ( .o(_net_10467), .ck(clk), .d(n1145) );
ms00f80  l0134 ( .o(_net_10417), .ck(clk), .d(n1150) );
ms00f80  l0135 ( .o(net_10530), .ck(clk), .d(n1155) );
ms00f80  l0136 ( .o(_net_9171), .ck(clk), .d(n1160) );
ms00f80  l0137 ( .o(net_9767), .ck(clk), .d(n1165) );
ms00f80  l0138 ( .o(_net_9375), .ck(clk), .d(n1170) );
ms00f80  l0139 ( .o(net_10518), .ck(clk), .d(n1175) );
ms00f80  l0140 ( .o(x589), .ck(clk), .d(n1179) );
ms00f80  l0141 ( .o(_net_9394), .ck(clk), .d(n1183) );
ms00f80  l0142 ( .o(_net_10411), .ck(clk), .d(n1188) );
ms00f80  l0143 ( .o(net_9274), .ck(clk), .d(n1193) );
ms00f80  l0144 ( .o(_net_10156), .ck(clk), .d(n1198) );
ms00f80  l0145 ( .o(net_9912), .ck(clk), .d(n1203) );
ms00f80  l0146 ( .o(net_9948), .ck(clk), .d(n1208) );
ms00f80  l0147 ( .o(_net_10368), .ck(clk), .d(n1213) );
ms00f80  l0148 ( .o(x1240), .ck(clk), .d(n1218) );
ms00f80  l0149 ( .o(net_9965), .ck(clk), .d(n1222) );
ms00f80  l0150 ( .o(net_10484), .ck(clk), .d(n1227) );
ms00f80  l0151 ( .o(_net_9751), .ck(clk), .d(n1232) );
ms00f80  l0152 ( .o(_net_10243), .ck(clk), .d(n1237) );
ms00f80  l0153 ( .o(_net_8833), .ck(clk), .d(n1242) );
ms00f80  l0154 ( .o(net_206), .ck(clk), .d(n1247) );
ms00f80  l0155 ( .o(net_10084), .ck(clk), .d(n1252) );
ms00f80  l0156 ( .o(net_9139), .ck(clk), .d(n1257) );
ms00f80  l0157 ( .o(_net_10319), .ck(clk), .d(n1262) );
ms00f80  l0158 ( .o(net_10181), .ck(clk), .d(n1267) );
ms00f80  l0159 ( .o(net_10021), .ck(clk), .d(n1272) );
ms00f80  l0160 ( .o(_net_163), .ck(clk), .d(n1277) );
ms00f80  l0161 ( .o(net_10303), .ck(clk), .d(n1282) );
ms00f80  l0162 ( .o(net_9859), .ck(clk), .d(n1286) );
ms00f80  l0163 ( .o(_net_10479), .ck(clk), .d(n1291) );
ms00f80  l0164 ( .o(_net_9552), .ck(clk), .d(n1296) );
ms00f80  l0165 ( .o(net_10059), .ck(clk), .d(n1301) );
ms00f80  l0166 ( .o(_net_9320), .ck(clk), .d(n1306) );
ms00f80  l0167 ( .o(net_9489), .ck(clk), .d(n1310) );
ms00f80  l0168 ( .o(net_9182), .ck(clk), .d(n1315) );
ms00f80  l0169 ( .o(_net_9932), .ck(clk), .d(n1320) );
ms00f80  l0170 ( .o(net_9902), .ck(clk), .d(n1325) );
ms00f80  l0171 ( .o(net_9860), .ck(clk), .d(n1330) );
ms00f80  l0172 ( .o(net_9454), .ck(clk), .d(n1335) );
ms00f80  l0173 ( .o(net_9978), .ck(clk), .d(n1339) );
ms00f80  l0174 ( .o(net_9924), .ck(clk), .d(n1344) );
ms00f80  l0175 ( .o(_net_155), .ck(clk), .d(n1349) );
ms00f80  l0176 ( .o(net_9127), .ck(clk), .d(n1354) );
ms00f80  l0177 ( .o(net_9677), .ck(clk), .d(n1359) );
ms00f80  l0178 ( .o(net_258), .ck(clk), .d(n1364) );
ms00f80  l0179 ( .o(_net_9177), .ck(clk), .d(n1369) );
ms00f80  l0180 ( .o(_net_158), .ck(clk), .d(n1374) );
ms00f80  l0181 ( .o(_net_10336), .ck(clk), .d(n1379) );
ms00f80  l0182 ( .o(_net_9536), .ck(clk), .d(n1384) );
ms00f80  l0183 ( .o(net_9281), .ck(clk), .d(n1388) );
ms00f80  l0184 ( .o(net_228), .ck(clk), .d(n1392) );
ms00f80  l0185 ( .o(net_9286), .ck(clk), .d(n1397) );
ms00f80  l0186 ( .o(_net_9649), .ck(clk), .d(n1401) );
ms00f80  l0187 ( .o(_net_10375), .ck(clk), .d(n1406) );
ms00f80  l0188 ( .o(x1121), .ck(clk), .d(n1411) );
ms00f80  l0189 ( .o(net_10180), .ck(clk), .d(n1415) );
ms00f80  l0190 ( .o(_net_10126), .ck(clk), .d(n1420) );
ms00f80  l0191 ( .o(_net_9930), .ck(clk), .d(n1425) );
ms00f80  l0192 ( .o(net_313), .ck(clk), .d(n1430) );
ms00f80  l0193 ( .o(net_9647), .ck(clk), .d(n1435) );
ms00f80  l0194 ( .o(net_299), .ck(clk), .d(n1440) );
ms00f80  l0195 ( .o(net_9665), .ck(clk), .d(n1444) );
ms00f80  l0196 ( .o(_net_9245), .ck(clk), .d(n1449) );
ms00f80  l0197 ( .o(net_9626), .ck(clk), .d(n1454) );
ms00f80  l0198 ( .o(_net_9590), .ck(clk), .d(n1459) );
ms00f80  l0199 ( .o(net_9815), .ck(clk), .d(n1464) );
ms00f80  l0200 ( .o(_net_10158), .ck(clk), .d(n1469) );
ms00f80  l0201 ( .o(x1113), .ck(clk), .d(n1474) );
ms00f80  l0202 ( .o(net_9218), .ck(clk), .d(n1478) );
ms00f80  l0203 ( .o(net_9814), .ck(clk), .d(n1483) );
ms00f80  l0204 ( .o(net_9338), .ck(clk), .d(n1488) );
ms00f80  l0205 ( .o(net_100), .ck(clk), .d(n1492) );
ms00f80  l0206 ( .o(_net_10061), .ck(clk), .d(n1497) );
ms00f80  l0207 ( .o(net_9848), .ck(clk), .d(n1502) );
ms00f80  l0208 ( .o(_net_8846), .ck(clk), .d(n1507) );
ms00f80  l0209 ( .o(_net_10366), .ck(clk), .d(n1512) );
ms00f80  l0210 ( .o(net_305), .ck(clk), .d(n1517) );
ms00f80  l0211 ( .o(_net_9186), .ck(clk), .d(n1521) );
ms00f80  l0212 ( .o(net_9722), .ck(clk), .d(n1526) );
ms00f80  l0213 ( .o(net_10193), .ck(clk), .d(n1531) );
ms00f80  l0214 ( .o(net_9330), .ck(clk), .d(n1536) );
ms00f80  l0215 ( .o(net_9856), .ck(clk), .d(n1540) );
ms00f80  l0216 ( .o(net_9456), .ck(clk), .d(n1545) );
ms00f80  l0217 ( .o(_net_10331), .ck(clk), .d(n1549) );
ms00f80  l0218 ( .o(net_9849), .ck(clk), .d(n1554) );
ms00f80  l0219 ( .o(net_9143), .ck(clk), .d(n1559) );
ms00f80  l0220 ( .o(net_9826), .ck(clk), .d(n1564) );
ms00f80  l0221 ( .o(net_9988), .ck(clk), .d(n1569) );
ms00f80  l0222 ( .o(net_10045), .ck(clk), .d(n1574) );
ms00f80  l0223 ( .o(x1197), .ck(clk), .d(n1579) );
ms00f80  l0224 ( .o(net_97), .ck(clk), .d(n1582) );
ms00f80  l0225 ( .o(net_9708), .ck(clk), .d(n1587) );
ms00f80  l0226 ( .o(_net_10113), .ck(clk), .d(n1592) );
ms00f80  l0227 ( .o(_net_10326), .ck(clk), .d(n1597) );
ms00f80  l0228 ( .o(net_311), .ck(clk), .d(n1602) );
ms00f80  l0229 ( .o(x1290), .ck(clk), .d(n1605) );
ms00f80  l0230 ( .o(net_10047), .ck(clk), .d(n1609) );
ms00f80  l0231 ( .o(_net_9313), .ck(clk), .d(n1614) );
ms00f80  l0232 ( .o(_net_9267), .ck(clk), .d(n1618) );
ms00f80  l0233 ( .o(net_9303), .ck(clk), .d(n1623) );
ms00f80  l0234 ( .o(net_302), .ck(clk), .d(n1627) );
ms00f80  l0235 ( .o(_net_10217), .ck(clk), .d(n1631) );
ms00f80  l0236 ( .o(_net_9322), .ck(clk), .d(n1636) );
ms00f80  l0237 ( .o(_net_9736), .ck(clk), .d(n1641) );
ms00f80  l0238 ( .o(net_9981), .ck(clk), .d(n1646) );
ms00f80  l0239 ( .o(net_10077), .ck(clk), .d(n1651) );
ms00f80  l0240 ( .o(net_9672), .ck(clk), .d(n1656) );
ms00f80  l0241 ( .o(_net_9512), .ck(clk), .d(n1661) );
ms00f80  l0242 ( .o(net_9577), .ck(clk), .d(n1666) );
ms00f80  l0243 ( .o(net_9367), .ck(clk), .d(n1671) );
ms00f80  l0244 ( .o(net_9954), .ck(clk), .d(n1676) );
ms00f80  l0245 ( .o(_net_9390), .ck(clk), .d(n1681) );
ms00f80  l0246 ( .o(_net_9302), .ck(clk), .d(n1686) );
ms00f80  l0247 ( .o(net_107), .ck(clk), .d(n1691) );
ms00f80  l0248 ( .o(net_9654), .ck(clk), .d(n1696) );
ms00f80  l0249 ( .o(_net_10307), .ck(clk), .d(n1701) );
ms00f80  l0250 ( .o(net_9350), .ck(clk), .d(n1706) );
ms00f80  l0251 ( .o(_net_9637), .ck(clk), .d(n1711) );
ms00f80  l0252 ( .o(net_9500), .ck(clk), .d(n1715) );
ms00f80  l0253 ( .o(net_10081), .ck(clk), .d(n1720) );
ms00f80  l0254 ( .o(_net_10440), .ck(clk), .d(n1725) );
ms00f80  l0255 ( .o(net_9893), .ck(clk), .d(n1730) );
ms00f80  l0256 ( .o(net_9451), .ck(clk), .d(n1735) );
ms00f80  l0257 ( .o(net_9695), .ck(clk), .d(n1739) );
ms00f80  l0258 ( .o(net_9801), .ck(clk), .d(n1744) );
ms00f80  l0259 ( .o(_net_9419), .ck(clk), .d(n1749) );
ms00f80  l0260 ( .o(_net_9827), .ck(clk), .d(n1754) );
ms00f80  l0261 ( .o(_net_9292), .ck(clk), .d(n1759) );
ms00f80  l0262 ( .o(net_10135), .ck(clk), .d(n1764) );
ms00f80  l0263 ( .o(net_10190), .ck(clk), .d(n1769) );
ms00f80  l0264 ( .o(net_9199), .ck(clk), .d(n1774) );
ms00f80  l0265 ( .o(net_9180), .ck(clk), .d(n1779) );
ms00f80  l0266 ( .o(net_92), .ck(clk), .d(n1783) );
ms00f80  l0267 ( .o(net_9951), .ck(clk), .d(n1787) );
ms00f80  l0268 ( .o(_net_9633), .ck(clk), .d(n1792) );
ms00f80  l0269 ( .o(_net_9424), .ck(clk), .d(n1797) );
ms00f80  l0270 ( .o(_net_9372), .ck(clk), .d(n1802) );
ms00f80  l0271 ( .o(net_9435), .ck(clk), .d(n1807) );
ms00f80  l0272 ( .o(_net_10115), .ck(clk), .d(n1812) );
ms00f80  l0273 ( .o(_net_9600), .ck(clk), .d(n1817) );
ms00f80  l0274 ( .o(_net_10347), .ck(clk), .d(n1822) );
ms00f80  l0275 ( .o(net_9479), .ck(clk), .d(n1826) );
ms00f80  l0276 ( .o(x1206), .ck(clk), .d(n1831) );
ms00f80  l0277 ( .o(_net_127), .ck(clk), .d(n1835) );
ms00f80  l0278 ( .o(net_9159), .ck(clk), .d(n1839) );
ms00f80  l0279 ( .o(_net_10271), .ck(clk), .d(n1844) );
ms00f80  l0280 ( .o(_net_10227), .ck(clk), .d(n1849) );
ms00f80  l0281 ( .o(_net_9317), .ck(clk), .d(n1854) );
ms00f80  l0282 ( .o(net_9738), .ck(clk), .d(n1859) );
ms00f80  l0283 ( .o(net_9473), .ck(clk), .d(n1863) );
ms00f80  l0284 ( .o(_net_157), .ck(clk), .d(n1868) );
ms00f80  l0285 ( .o(net_9481), .ck(clk), .d(n1872) );
ms00f80  l0286 ( .o(net_10020), .ck(clk), .d(n1877) );
ms00f80  l0287 ( .o(_net_9191), .ck(clk), .d(n1881) );
ms00f80  l0288 ( .o(_net_10511), .ck(clk), .d(n1886) );
ms00f80  l0289 ( .o(net_10239), .ck(clk), .d(n1891) );
ms00f80  l0290 ( .o(_net_10359), .ck(clk), .d(n1896) );
ms00f80  l0291 ( .o(_net_268), .ck(clk), .d(n1901) );
ms00f80  l0292 ( .o(net_9576), .ck(clk), .d(n1906) );
ms00f80  l0293 ( .o(_net_265), .ck(clk), .d(n1911) );
ms00f80  l0294 ( .o(_net_9380), .ck(clk), .d(n1916) );
ms00f80  l0295 ( .o(net_10497), .ck(clk), .d(n1921) );
ms00f80  l0296 ( .o(_net_187), .ck(clk), .d(n1926) );
ms00f80  l0297 ( .o(net_9347), .ck(clk), .d(n1931) );
ms00f80  l0298 ( .o(_net_8817), .ck(clk), .d(n1936) );
ms00f80  l0299 ( .o(_net_10231), .ck(clk), .d(n1941) );
ms00f80  l0300 ( .o(net_10493), .ck(clk), .d(n1946) );
ms00f80  l0301 ( .o(_net_10420), .ck(clk), .d(n1951) );
ms00f80  l0302 ( .o(net_9137), .ck(clk), .d(n1956) );
ms00f80  l0303 ( .o(net_10178), .ck(clk), .d(n1960) );
ms00f80  l0304 ( .o(_net_10369), .ck(clk), .d(n1965) );
ms00f80  l0305 ( .o(net_9684), .ck(clk), .d(n1970) );
ms00f80  l0306 ( .o(net_9578), .ck(clk), .d(n1975) );
ms00f80  l0307 ( .o(net_9614), .ck(clk), .d(n1980) );
ms00f80  l0308 ( .o(_net_10091), .ck(clk), .d(n1985) );
ms00f80  l0309 ( .o(net_9891), .ck(clk), .d(n1990) );
ms00f80  l0310 ( .o(net_9998), .ck(clk), .d(n1995) );
ms00f80  l0311 ( .o(_net_10487), .ck(clk), .d(n2000) );
ms00f80  l0312 ( .o(net_9808), .ck(clk), .d(n2005) );
ms00f80  l0313 ( .o(net_9996), .ck(clk), .d(n2010) );
ms00f80  l0314 ( .o(_net_10452), .ck(clk), .d(n2015) );
ms00f80  l0315 ( .o(_net_10373), .ck(clk), .d(n2020) );
ms00f80  l0316 ( .o(_net_10252), .ck(clk), .d(n2025) );
ms00f80  l0317 ( .o(net_10290), .ck(clk), .d(n2030) );
ms00f80  l0318 ( .o(_net_10443), .ck(clk), .d(n2035) );
ms00f80  l0319 ( .o(net_8818), .ck(clk), .d(n2040) );
ms00f80  l0320 ( .o(_net_9318), .ck(clk), .d(n2045) );
ms00f80  l0321 ( .o(_net_9850), .ck(clk), .d(n2050) );
ms00f80  l0322 ( .o(net_9901), .ck(clk), .d(n2055) );
ms00f80  l0323 ( .o(_net_8828), .ck(clk), .d(n2060) );
ms00f80  l0324 ( .o(_net_202), .ck(clk), .d(n2065) );
ms00f80  l0325 ( .o(_net_10090), .ck(clk), .d(n2070) );
ms00f80  l0326 ( .o(_net_9213), .ck(clk), .d(n2075) );
ms00f80  l0327 ( .o(_net_9396), .ck(clk), .d(n2080) );
ms00f80  l0328 ( .o(_net_10528), .ck(clk), .d(n2085) );
ms00f80  l0329 ( .o(_net_9563), .ck(clk), .d(n2090) );
ms00f80  l0330 ( .o(_net_10224), .ck(clk), .d(n2095) );
ms00f80  l0331 ( .o(_net_10123), .ck(clk), .d(n2100) );
ms00f80  l0332 ( .o(_net_10435), .ck(clk), .d(n2105) );
ms00f80  l0333 ( .o(_net_10103), .ck(clk), .d(n2110) );
ms00f80  l0334 ( .o(_net_10098), .ck(clk), .d(n2115) );
ms00f80  l0335 ( .o(_net_10262), .ck(clk), .d(n2120) );
ms00f80  l0336 ( .o(net_208), .ck(clk), .d(n2125) );
ms00f80  l0337 ( .o(_net_10446), .ck(clk), .d(n2130) );
ms00f80  l0338 ( .o(net_9528), .ck(clk), .d(n2135) );
ms00f80  l0339 ( .o(_net_9351), .ck(clk), .d(n2140) );
ms00f80  l0340 ( .o(net_9761), .ck(clk), .d(n2145) );
ms00f80  l0341 ( .o(net_9972), .ck(clk), .d(n2150) );
ms00f80  l0342 ( .o(net_9894), .ck(clk), .d(n2155) );
ms00f80  l0343 ( .o(_net_10543), .ck(clk), .d(n2160) );
ms00f80  l0344 ( .o(_net_9639), .ck(clk), .d(n2165) );
ms00f80  l0345 ( .o(net_9158), .ck(clk), .d(n2169) );
ms00f80  l0346 ( .o(_net_10483), .ck(clk), .d(n2174) );
ms00f80  l0347 ( .o(net_9913), .ck(clk), .d(n2179) );
ms00f80  l0348 ( .o(_net_125), .ck(clk), .d(n2184) );
ms00f80  l0349 ( .o(x1129), .ck(clk), .d(n2189) );
ms00f80  l0350 ( .o(net_10039), .ck(clk), .d(n2193) );
ms00f80  l0351 ( .o(net_214), .ck(clk), .d(n2198) );
ms00f80  l0352 ( .o(net_10409), .ck(clk), .d(n2202) );
ms00f80  l0353 ( .o(net_9579), .ck(clk), .d(n2207) );
ms00f80  l0354 ( .o(_net_10311), .ck(clk), .d(n2212) );
ms00f80  l0355 ( .o(net_256), .ck(clk), .d(n2217) );
ms00f80  l0356 ( .o(net_10050), .ck(clk), .d(n2222) );
ms00f80  l0357 ( .o(_net_9437), .ck(clk), .d(n2227) );
ms00f80  l0358 ( .o(_net_10413), .ck(clk), .d(n2232) );
ms00f80  l0359 ( .o(net_213), .ck(clk), .d(n2237) );
ms00f80  l0360 ( .o(_net_9640), .ck(clk), .d(n2242) );
ms00f80  l0361 ( .o(net_10093), .ck(clk), .d(n2246) );
ms00f80  l0362 ( .o(_net_10357), .ck(clk), .d(n2251) );
ms00f80  l0363 ( .o(net_9527), .ck(clk), .d(n2256) );
ms00f80  l0364 ( .o(net_9878), .ck(clk), .d(n2261) );
ms00f80  l0365 ( .o(net_215), .ck(clk), .d(n2266) );
ms00f80  l0366 ( .o(_net_10382), .ck(clk), .d(n2271) );
ms00f80  l0367 ( .o(_net_10226), .ck(clk), .d(n2276) );
ms00f80  l0368 ( .o(net_9962), .ck(clk), .d(n2281) );
ms00f80  l0369 ( .o(net_9883), .ck(clk), .d(n2286) );
ms00f80  l0370 ( .o(net_9544), .ck(clk), .d(n2291) );
ms00f80  l0371 ( .o(net_9710), .ck(clk), .d(n2296) );
ms00f80  l0372 ( .o(net_10194), .ck(clk), .d(n2301) );
ms00f80  l0373 ( .o(net_9653), .ck(clk), .d(n2306) );
ms00f80  l0374 ( .o(_net_10468), .ck(clk), .d(n2311) );
ms00f80  l0375 ( .o(net_9794), .ck(clk), .d(n2316) );
ms00f80  l0376 ( .o(net_9525), .ck(clk), .d(n2321) );
ms00f80  l0377 ( .o(net_90), .ck(clk), .d(n2325) );
ms00f80  l0378 ( .o(net_9116), .ck(clk), .d(n2330) );
ms00f80  l0379 ( .o(x1223), .ck(clk), .d(n2334) );
ms00f80  l0380 ( .o(net_282), .ck(clk), .d(n2338) );
ms00f80  l0381 ( .o(net_149), .ck(clk), .d(n2342) );
ms00f80  l0382 ( .o(net_9151), .ck(clk), .d(n2347) );
ms00f80  l0383 ( .o(_net_10371), .ck(clk), .d(n2352) );
ms00f80  l0384 ( .o(net_9679), .ck(clk), .d(n2357) );
ms00f80  l0385 ( .o(net_9900), .ck(clk), .d(n2362) );
ms00f80  l0386 ( .o(net_9253), .ck(clk), .d(n2367) );
ms00f80  l0387 ( .o(x555), .ck(clk), .d(n2371) );
ms00f80  l0388 ( .o(_net_130), .ck(clk), .d(n2375) );
ms00f80  l0389 ( .o(_net_9938), .ck(clk), .d(n2380) );
ms00f80  l0390 ( .o(_net_10174), .ck(clk), .d(n2385) );
ms00f80  l0391 ( .o(net_10508), .ck(clk), .d(n2390) );
ms00f80  l0392 ( .o(net_9585), .ck(clk), .d(n2395) );
ms00f80  l0393 ( .o(net_9750), .ck(clk), .d(n2400) );
ms00f80  l0394 ( .o(net_9360), .ck(clk), .d(n2404) );
ms00f80  l0395 ( .o(_net_10489), .ck(clk), .d(n2409) );
ms00f80  l0396 ( .o(_net_9660), .ck(clk), .d(n2414) );
ms00f80  l0397 ( .o(net_10176), .ck(clk), .d(n2419) );
ms00f80  l0398 ( .o(_net_10461), .ck(clk), .d(n2424) );
ms00f80  l0399 ( .o(_net_9185), .ck(clk), .d(n2429) );
ms00f80  l0400 ( .o(_net_10127), .ck(clk), .d(n2434) );
ms00f80  l0401 ( .o(net_9610), .ck(clk), .d(n2439) );
ms00f80  l0402 ( .o(_net_9835), .ck(clk), .d(n2444) );
ms00f80  l0403 ( .o(net_9256), .ck(clk), .d(n2449) );
ms00f80  l0404 ( .o(net_9487), .ck(clk), .d(n2453) );
ms00f80  l0405 ( .o(_net_259), .ck(clk), .d(n2458) );
ms00f80  l0406 ( .o(net_10506), .ck(clk), .d(n2463) );
ms00f80  l0407 ( .o(net_9181), .ck(clk), .d(n2468) );
ms00f80  l0408 ( .o(net_9305), .ck(clk), .d(n2473) );
ms00f80  l0409 ( .o(net_9205), .ck(clk), .d(n2477) );
ms00f80  l0410 ( .o(_net_9354), .ck(clk), .d(n2482) );
ms00f80  l0411 ( .o(_net_10374), .ck(clk), .d(n2487) );
ms00f80  l0412 ( .o(net_9947), .ck(clk), .d(n2492) );
ms00f80  l0413 ( .o(_net_9193), .ck(clk), .d(n2497) );
ms00f80  l0414 ( .o(_net_9642), .ck(clk), .d(n2502) );
ms00f80  l0415 ( .o(net_10192), .ck(clk), .d(n2507) );
ms00f80  l0416 ( .o(net_264), .ck(clk), .d(n2512) );
ms00f80  l0417 ( .o(_net_8829), .ck(clk), .d(n2517) );
ms00f80  l0418 ( .o(_net_9300), .ck(clk), .d(n2522) );
ms00f80  l0419 ( .o(net_9846), .ck(clk), .d(n2527) );
ms00f80  l0420 ( .o(net_10526), .ck(clk), .d(n2532) );
ms00f80  l0421 ( .o(net_9452), .ck(clk), .d(n2537) );
ms00f80  l0422 ( .o(_net_10351), .ck(clk), .d(n2541) );
ms00f80  l0423 ( .o(net_9570), .ck(clk), .d(n2546) );
ms00f80  l0424 ( .o(_net_9927), .ck(clk), .d(n2551) );
ms00f80  l0425 ( .o(net_140), .ck(clk), .d(n2556) );
ms00f80  l0426 ( .o(x480), .ck(clk), .d(n2560) );
ms00f80  l0427 ( .o(net_9652), .ck(clk), .d(n2564) );
ms00f80  l0428 ( .o(x798), .ck(clk), .d(n2568) );
ms00f80  l0429 ( .o(net_10240), .ck(clk), .d(n2572) );
ms00f80  l0430 ( .o(net_10008), .ck(clk), .d(n2577) );
ms00f80  l0431 ( .o(_net_10318), .ck(clk), .d(n2582) );
ms00f80  l0432 ( .o(net_9224), .ck(clk), .d(n2587) );
ms00f80  l0433 ( .o(net_9788), .ck(clk), .d(n2592) );
ms00f80  l0434 ( .o(_net_10363), .ck(clk), .d(n2597) );
ms00f80  l0435 ( .o(net_9960), .ck(clk), .d(n2602) );
ms00f80  l0436 ( .o(_net_10349), .ck(clk), .d(n2607) );
ms00f80  l0437 ( .o(_net_10384), .ck(clk), .d(n2612) );
ms00f80  l0438 ( .o(_net_165), .ck(clk), .d(n2617) );
ms00f80  l0439 ( .o(net_9540), .ck(clk), .d(n2622) );
ms00f80  l0440 ( .o(net_10058), .ck(clk), .d(n2627) );
ms00f80  l0441 ( .o(_net_270), .ck(clk), .d(n2632) );
ms00f80  l0442 ( .o(net_9228), .ck(clk), .d(n2637) );
ms00f80  l0443 ( .o(_net_184), .ck(clk), .d(n2642) );
ms00f80  l0444 ( .o(net_10536), .ck(clk), .d(n2647) );
ms00f80  l0445 ( .o(_net_10101), .ck(clk), .d(n2652) );
ms00f80  l0446 ( .o(_net_183), .ck(clk), .d(n2657) );
ms00f80  l0447 ( .o(_net_9561), .ck(clk), .d(n2662) );
ms00f80  l0448 ( .o(net_9132), .ck(clk), .d(n2667) );
ms00f80  l0449 ( .o(net_9898), .ck(clk), .d(n2671) );
ms00f80  l0450 ( .o(_net_267), .ck(clk), .d(n2676) );
ms00f80  l0451 ( .o(net_10380), .ck(clk), .d(n2681) );
ms00f80  l0452 ( .o(net_196), .ck(clk), .d(n2685) );
ms00f80  l0453 ( .o(net_9634), .ck(clk), .d(n2690) );
ms00f80  l0454 ( .o(net_9275), .ck(clk), .d(n2695) );
ms00f80  l0455 ( .o(_net_10352), .ck(clk), .d(n2700) );
ms00f80  l0456 ( .o(net_9220), .ck(clk), .d(n2705) );
ms00f80  l0457 ( .o(net_145), .ck(clk), .d(n2710) );
ms00f80  l0458 ( .o(net_10494), .ck(clk), .d(n2715) );
ms00f80  l0459 ( .o(net_10539), .ck(clk), .d(n2720) );
ms00f80  l0460 ( .o(net_10011), .ck(clk), .d(n2725) );
ms00f80  l0461 ( .o(_net_8844), .ck(clk), .d(n2730) );
ms00f80  l0462 ( .o(_net_117), .ck(clk), .d(n2735) );
ms00f80  l0463 ( .o(net_9607), .ck(clk), .d(n2740) );
ms00f80  l0464 ( .o(_net_191), .ck(clk), .d(n2745) );
ms00f80  l0465 ( .o(_net_9420), .ck(clk), .d(n2750) );
ms00f80  l0466 ( .o(_net_10436), .ck(clk), .d(n2755) );
ms00f80  l0467 ( .o(_net_10048), .ck(clk), .d(n2760) );
ms00f80  l0468 ( .o(_net_9383), .ck(clk), .d(n2765) );
ms00f80  l0469 ( .o(net_9493), .ck(clk), .d(n2769) );
ms00f80  l0470 ( .o(_net_9201), .ck(clk), .d(n2774) );
ms00f80  l0471 ( .o(_net_9745), .ck(clk), .d(n2779) );
ms00f80  l0472 ( .o(_net_10031), .ck(clk), .d(n2784) );
ms00f80  l0473 ( .o(_net_9241), .ck(clk), .d(n2789) );
ms00f80  l0474 ( .o(net_10490), .ck(clk), .d(n2794) );
ms00f80  l0475 ( .o(net_9483), .ck(clk), .d(n2798) );
ms00f80  l0476 ( .o(net_106), .ck(clk), .d(n2803) );
ms00f80  l0477 ( .o(net_103), .ck(clk), .d(n2808) );
ms00f80  l0478 ( .o(net_9881), .ck(clk), .d(n2813) );
ms00f80  l0479 ( .o(net_9495), .ck(clk), .d(n2817) );
ms00f80  l0480 ( .o(net_10507), .ck(clk), .d(n2822) );
ms00f80  l0481 ( .o(_net_9573), .ck(clk), .d(n2827) );
ms00f80  l0482 ( .o(net_9438), .ck(clk), .d(n2832) );
ms00f80  l0483 ( .o(_net_9246), .ck(clk), .d(n2836) );
ms00f80  l0484 ( .o(net_9802), .ck(clk), .d(n2841) );
ms00f80  l0485 ( .o(_net_9236), .ck(clk), .d(n2846) );
ms00f80  l0486 ( .o(net_9333), .ck(clk), .d(n2851) );
ms00f80  l0487 ( .o(net_10072), .ck(clk), .d(n2855) );
ms00f80  l0488 ( .o(x494), .ck(clk), .d(n2860) );
ms00f80  l0489 ( .o(net_10295), .ck(clk), .d(n2864) );
ms00f80  l0490 ( .o(_net_10361), .ck(clk), .d(n2869) );
ms00f80  l0491 ( .o(x747), .ck(clk), .d(n2874) );
ms00f80  l0492 ( .o(_net_181), .ck(clk), .d(n2878) );
ms00f80  l0493 ( .o(_net_9744), .ck(clk), .d(n2883) );
ms00f80  l0494 ( .o(net_9905), .ck(clk), .d(n2888) );
ms00f80  l0495 ( .o(_net_10253), .ck(clk), .d(n2893) );
ms00f80  l0496 ( .o(net_10448), .ck(clk), .d(n2898) );
ms00f80  l0497 ( .o(net_9575), .ck(clk), .d(n2903) );
ms00f80  l0498 ( .o(net_9439), .ck(clk), .d(n2908) );
ms00f80  l0499 ( .o(_net_9404), .ck(clk), .d(n2912) );
ms00f80  l0500 ( .o(net_10393), .ck(clk), .d(n2917) );
ms00f80  l0501 ( .o(net_9908), .ck(clk), .d(n2922) );
ms00f80  l0502 ( .o(_net_9190), .ck(clk), .d(n2927) );
ms00f80  l0503 ( .o(net_10002), .ck(clk), .d(n2932) );
ms00f80  l0504 ( .o(_net_10033), .ck(clk), .d(n2937) );
ms00f80  l0505 ( .o(net_9441), .ck(clk), .d(n2942) );
ms00f80  l0506 ( .o(net_8836), .ck(clk), .d(n2946) );
ms00f80  l0507 ( .o(_net_9580), .ck(clk), .d(n2951) );
ms00f80  l0508 ( .o(x447), .ck(clk), .d(n2956) );
ms00f80  l0509 ( .o(_net_9828), .ck(clk), .d(n2960) );
ms00f80  l0510 ( .o(_net_9377), .ck(clk), .d(n2965) );
ms00f80  l0511 ( .o(_net_9417), .ck(clk), .d(n2970) );
ms00f80  l0512 ( .o(_net_9731), .ck(clk), .d(n2975) );
ms00f80  l0513 ( .o(_net_10335), .ck(clk), .d(n2980) );
ms00f80  l0514 ( .o(net_211), .ck(clk), .d(n2985) );
ms00f80  l0515 ( .o(_net_10206), .ck(clk), .d(n2990) );
ms00f80  l0516 ( .o(net_9952), .ck(clk), .d(n2995) );
ms00f80  l0517 ( .o(net_9984), .ck(clk), .d(n3000) );
ms00f80  l0518 ( .o(_net_124), .ck(clk), .d(n3005) );
ms00f80  l0519 ( .o(_net_10054), .ck(clk), .d(n3010) );
ms00f80  l0520 ( .o(net_9970), .ck(clk), .d(n3015) );
ms00f80  l0521 ( .o(_net_9062), .ck(clk), .d(n3020) );
ms00f80  l0522 ( .o(_net_9370), .ck(clk), .d(n3025) );
ms00f80  l0523 ( .o(_net_10333), .ck(clk), .d(n3030) );
ms00f80  l0524 ( .o(net_9496), .ck(clk), .d(n3034) );
ms00f80  l0525 ( .o(x465), .ck(clk), .d(n3039) );
ms00f80  l0526 ( .o(_net_10451), .ck(clk), .d(n3043) );
ms00f80  l0527 ( .o(_net_9314), .ck(clk), .d(n3048) );
ms00f80  l0528 ( .o(_net_10414), .ck(clk), .d(n3053) );
ms00f80  l0529 ( .o(net_9533), .ck(clk), .d(n3058) );
ms00f80  l0530 ( .o(net_221), .ck(clk), .d(n3063) );
ms00f80  l0531 ( .o(_net_10163), .ck(clk), .d(n3068) );
ms00f80  l0532 ( .o(net_285), .ck(clk), .d(n3073) );
ms00f80  l0533 ( .o(_net_10362), .ck(clk), .d(n3077) );
ms00f80  l0534 ( .o(net_9816), .ck(clk), .d(n3082) );
ms00f80  l0535 ( .o(_net_10309), .ck(clk), .d(n3087) );
ms00f80  l0536 ( .o(_net_10107), .ck(clk), .d(n3092) );
ms00f80  l0537 ( .o(net_296), .ck(clk), .d(n3097) );
ms00f80  l0538 ( .o(net_9673), .ck(clk), .d(n3101) );
ms00f80  l0539 ( .o(net_9162), .ck(clk), .d(n3106) );
ms00f80  l0540 ( .o(_net_9167), .ck(clk), .d(n3111) );
ms00f80  l0541 ( .o(_net_9294), .ck(clk), .d(n3116) );
ms00f80  l0542 ( .o(net_9650), .ck(clk), .d(n3121) );
ms00f80  l0543 ( .o(_net_9323), .ck(clk), .d(n3126) );
ms00f80  l0544 ( .o(net_9273), .ck(clk), .d(n3131) );
ms00f80  l0545 ( .o(_net_10025), .ck(clk), .d(n3136) );
ms00f80  l0546 ( .o(net_10175), .ck(clk), .d(n3141) );
ms00f80  l0547 ( .o(_net_8845), .ck(clk), .d(n3146) );
ms00f80  l0548 ( .o(_net_9298), .ck(clk), .d(n3151) );
ms00f80  l0549 ( .o(net_9723), .ck(clk), .d(n3156) );
ms00f80  l0550 ( .o(net_9255), .ck(clk), .d(n3161) );
ms00f80  l0551 ( .o(net_9963), .ck(clk), .d(n3166) );
ms00f80  l0552 ( .o(_net_10129), .ck(clk), .d(n3171) );
ms00f80  l0553 ( .o(_net_152), .ck(clk), .d(n3176) );
ms00f80  l0554 ( .o(net_10068), .ck(clk), .d(n3181) );
ms00f80  l0555 ( .o(_net_9319), .ck(clk), .d(n3186) );
ms00f80  l0556 ( .o(net_9582), .ck(clk), .d(n3191) );
ms00f80  l0557 ( .o(net_9773), .ck(clk), .d(n3195) );
ms00f80  l0558 ( .o(net_10189), .ck(clk), .d(n3200) );
ms00f80  l0559 ( .o(net_9804), .ck(clk), .d(n3205) );
ms00f80  l0560 ( .o(net_9265), .ck(clk), .d(n3210) );
ms00f80  l0561 ( .o(net_9819), .ck(clk), .d(n3215) );
ms00f80  l0562 ( .o(net_9234), .ck(clk), .d(n3220) );
ms00f80  l0563 ( .o(net_9226), .ck(clk), .d(n3225) );
ms00f80  l0564 ( .o(net_9915), .ck(clk), .d(n3230) );
ms00f80  l0565 ( .o(x1357), .ck(clk), .d(n3234) );
ms00f80  l0566 ( .o(net_9886), .ck(clk), .d(n3238) );
ms00f80  l0567 ( .o(net_10073), .ck(clk), .d(n3243) );
ms00f80  l0568 ( .o(net_9492), .ck(clk), .d(n3247) );
ms00f80  l0569 ( .o(net_9656), .ck(clk), .d(n3252) );
ms00f80  l0570 ( .o(_net_9606), .ck(clk), .d(n3257) );
ms00f80  l0571 ( .o(_net_9183), .ck(clk), .d(n3262) );
ms00f80  l0572 ( .o(net_9922), .ck(clk), .d(n3267) );
ms00f80  l0573 ( .o(_net_9194), .ck(clk), .d(n3272) );
ms00f80  l0574 ( .o(net_244), .ck(clk), .d(n3277) );
ms00f80  l0575 ( .o(_net_10247), .ck(clk), .d(n3282) );
ms00f80  l0576 ( .o(net_101), .ck(clk), .d(n3287) );
ms00f80  l0577 ( .o(net_9155), .ck(clk), .d(n3291) );
ms00f80  l0578 ( .o(net_9184), .ck(clk), .d(n3296) );
ms00f80  l0579 ( .o(_net_9530), .ck(clk), .d(n3300) );
ms00f80  l0580 ( .o(_net_10229), .ck(clk), .d(n3305) );
ms00f80  l0581 ( .o(net_9359), .ck(clk), .d(n3310) );
ms00f80  l0582 ( .o(net_10296), .ck(clk), .d(n3315) );
ms00f80  l0583 ( .o(_net_9743), .ck(clk), .d(n3320) );
ms00f80  l0584 ( .o(net_9911), .ck(clk), .d(n3325) );
ms00f80  l0585 ( .o(net_10275), .ck(clk), .d(n3330) );
ms00f80  l0586 ( .o(_net_9242), .ck(clk), .d(n3335) );
ms00f80  l0587 ( .o(net_10291), .ck(clk), .d(n3340) );
ms00f80  l0588 ( .o(net_9792), .ck(clk), .d(n3345) );
ms00f80  l0589 ( .o(net_9680), .ck(clk), .d(n3350) );
ms00f80  l0590 ( .o(_net_10531), .ck(clk), .d(n3355) );
ms00f80  l0591 ( .o(net_250), .ck(clk), .d(n3359) );
ms00f80  l0592 ( .o(net_9625), .ck(clk), .d(n3364) );
ms00f80  l0593 ( .o(net_10503), .ck(clk), .d(n3369) );
ms00f80  l0594 ( .o(_net_10488), .ck(clk), .d(n3374) );
ms00f80  l0595 ( .o(net_9364), .ck(clk), .d(n3379) );
ms00f80  l0596 ( .o(_net_9434), .ck(clk), .d(n3384) );
ms00f80  l0597 ( .o(net_10533), .ck(clk), .d(n3389) );
ms00f80  l0598 ( .o(_net_9943), .ck(clk), .d(n3394) );
ms00f80  l0599 ( .o(net_10038), .ck(clk), .d(n3399) );
ms00f80  l0600 ( .o(_net_10434), .ck(clk), .d(n3404) );
ms00f80  l0601 ( .o(x1058), .ck(clk), .d(n3409) );
ms00f80  l0602 ( .o(net_9459), .ck(clk), .d(n3413) );
ms00f80  l0603 ( .o(net_249), .ck(clk), .d(n3416) );
ms00f80  l0604 ( .o(_net_10100), .ck(clk), .d(n3421) );
ms00f80  l0605 ( .o(net_9446), .ck(clk), .d(n3426) );
ms00f80  l0606 ( .o(net_10392), .ck(clk), .d(n3430) );
ms00f80  l0607 ( .o(net_210), .ck(clk), .d(n3435) );
ms00f80  l0608 ( .o(_net_10453), .ck(clk), .d(n3440) );
ms00f80  l0609 ( .o(net_9524), .ck(clk), .d(n3445) );
ms00f80  l0610 ( .o(net_9916), .ck(clk), .d(n3450) );
ms00f80  l0611 ( .o(_net_9608), .ck(clk), .d(n3455) );
ms00f80  l0612 ( .o(_net_10378), .ck(clk), .d(n3460) );
ms00f80  l0613 ( .o(_net_8843), .ck(clk), .d(n3465) );
ms00f80  l0614 ( .o(net_9786), .ck(clk), .d(n3470) );
ms00f80  l0615 ( .o(net_10387), .ck(clk), .d(n3475) );
ms00f80  l0616 ( .o(_net_8841), .ck(clk), .d(n3480) );
ms00f80  l0617 ( .o(net_10499), .ck(clk), .d(n3485) );
ms00f80  l0618 ( .o(_net_9601), .ck(clk), .d(n3490) );
ms00f80  l0619 ( .o(x1179), .ck(clk), .d(n3495) );
ms00f80  l0620 ( .o(net_262), .ck(clk), .d(n3499) );
ms00f80  l0621 ( .o(_net_9844), .ck(clk), .d(n3504) );
ms00f80  l0622 ( .o(x1095), .ck(clk), .d(n3509) );
ms00f80  l0623 ( .o(net_10009), .ck(clk), .d(n3513) );
ms00f80  l0624 ( .o(net_9782), .ck(clk), .d(n3518) );
ms00f80  l0625 ( .o(net_9212), .ck(clk), .d(n3523) );
ms00f80  l0626 ( .o(net_10496), .ck(clk), .d(n3528) );
ms00f80  l0627 ( .o(net_9522), .ck(clk), .d(n3533) );
ms00f80  l0628 ( .o(net_9785), .ck(clk), .d(n3538) );
ms00f80  l0629 ( .o(_net_10218), .ck(clk), .d(n3543) );
ms00f80  l0630 ( .o(_net_9172), .ck(clk), .d(n3548) );
ms00f80  l0631 ( .o(net_10195), .ck(clk), .d(n3553) );
ms00f80  l0632 ( .o(net_10394), .ck(clk), .d(n3558) );
ms00f80  l0633 ( .o(_net_9641), .ck(clk), .d(n3563) );
ms00f80  l0634 ( .o(_net_10225), .ck(clk), .d(n3568) );
ms00f80  l0635 ( .o(net_10284), .ck(clk), .d(n3573) );
ms00f80  l0636 ( .o(_net_10125), .ck(clk), .d(n3578) );
ms00f80  l0637 ( .o(_net_10220), .ck(clk), .d(n3583) );
ms00f80  l0638 ( .o(net_10294), .ck(clk), .d(n3588) );
ms00f80  l0639 ( .o(_net_172), .ck(clk), .d(n3593) );
ms00f80  l0640 ( .o(_net_10096), .ck(clk), .d(n3598) );
ms00f80  l0641 ( .o(net_10060), .ck(clk), .d(n3603) );
ms00f80  l0642 ( .o(net_9688), .ck(clk), .d(n3608) );
ms00f80  l0643 ( .o(net_10501), .ck(clk), .d(n3613) );
ms00f80  l0644 ( .o(net_218), .ck(clk), .d(n3618) );
ms00f80  l0645 ( .o(_net_9553), .ck(clk), .d(n3623) );
ms00f80  l0646 ( .o(net_9592), .ck(clk), .d(n3628) );
ms00f80  l0647 ( .o(net_9560), .ck(clk), .d(n3633) );
ms00f80  l0648 ( .o(x715), .ck(clk), .d(n3638) );
ms00f80  l0649 ( .o(net_10086), .ck(clk), .d(n3642) );
ms00f80  l0650 ( .o(_net_10512), .ck(clk), .d(n3647) );
ms00f80  l0651 ( .o(_net_10313), .ck(clk), .d(n3652) );
ms00f80  l0652 ( .o(net_9142), .ck(clk), .d(n3657) );
ms00f80  l0653 ( .o(_net_8824), .ck(clk), .d(n3662) );
ms00f80  l0654 ( .o(net_10016), .ck(clk), .d(n3667) );
ms00f80  l0655 ( .o(net_9775), .ck(clk), .d(n3672) );
ms00f80  l0656 ( .o(net_9769), .ck(clk), .d(n3677) );
ms00f80  l0657 ( .o(_net_10273), .ck(clk), .d(n3682) );
ms00f80  l0658 ( .o(_net_10473), .ck(clk), .d(n3687) );
ms00f80  l0659 ( .o(_net_10482), .ck(clk), .d(n3692) );
ms00f80  l0660 ( .o(net_9937), .ck(clk), .d(n3697) );
ms00f80  l0661 ( .o(_net_10209), .ck(clk), .d(n3702) );
ms00f80  l0662 ( .o(_net_10210), .ck(clk), .d(n3707) );
ms00f80  l0663 ( .o(_net_9385), .ck(clk), .d(n3712) );
ms00f80  l0664 ( .o(_net_9562), .ck(clk), .d(n3717) );
ms00f80  l0665 ( .o(_net_10372), .ck(clk), .d(n3722) );
ms00f80  l0666 ( .o(net_9811), .ck(clk), .d(n3727) );
ms00f80  l0667 ( .o(net_9862), .ck(clk), .d(n3732) );
ms00f80  l0668 ( .o(net_9523), .ck(clk), .d(n3737) );
ms00f80  l0669 ( .o(_net_9386), .ck(clk), .d(n3742) );
ms00f80  l0670 ( .o(net_10519), .ck(clk), .d(n3746) );
ms00f80  l0671 ( .o(_net_9829), .ck(clk), .d(n3750) );
ms00f80  l0672 ( .o(net_9471), .ck(clk), .d(n3754) );
ms00f80  l0673 ( .o(_net_9195), .ck(clk), .d(n3758) );
ms00f80  l0674 ( .o(net_109), .ck(clk), .d(n3763) );
ms00f80  l0675 ( .o(net_104), .ck(clk), .d(n3768) );
ms00f80  l0676 ( .o(_net_10242), .ck(clk), .d(n3773) );
ms00f80  l0677 ( .o(_net_10040), .ck(clk), .d(n3778) );
ms00f80  l0678 ( .o(net_99), .ck(clk), .d(n3782) );
ms00f80  l0679 ( .o(net_10132), .ck(clk), .d(n3787) );
ms00f80  l0680 ( .o(net_9468), .ck(clk), .d(n3792) );
ms00f80  l0681 ( .o(_net_10149), .ck(clk), .d(n3796) );
ms00f80  l0682 ( .o(x682), .ck(clk), .d(n3801) );
ms00f80  l0683 ( .o(net_9888), .ck(clk), .d(n3805) );
ms00f80  l0684 ( .o(net_10390), .ck(clk), .d(n3810) );
ms00f80  l0685 ( .o(net_9227), .ck(clk), .d(n3815) );
ms00f80  l0686 ( .o(_net_8823), .ck(clk), .d(n3820) );
ms00f80  l0687 ( .o(_net_9933), .ck(clk), .d(n3825) );
ms00f80  l0688 ( .o(_net_9344), .ck(clk), .d(n3830) );
ms00f80  l0689 ( .o(net_309), .ck(clk), .d(n3835) );
ms00f80  l0690 ( .o(net_9691), .ck(clk), .d(n3839) );
ms00f80  l0691 ( .o(net_9387), .ck(clk), .d(n3844) );
ms00f80  l0692 ( .o(net_9879), .ck(clk), .d(n3849) );
ms00f80  l0693 ( .o(_net_10328), .ck(clk), .d(n3854) );
ms00f80  l0694 ( .o(_net_275), .ck(clk), .d(n3859) );
ms00f80  l0695 ( .o(net_10001), .ck(clk), .d(n3864) );
ms00f80  l0696 ( .o(_net_274), .ck(clk), .d(n3869) );
ms00f80  l0697 ( .o(net_9230), .ck(clk), .d(n3874) );
ms00f80  l0698 ( .o(_net_10410), .ck(clk), .d(n3879) );
ms00f80  l0699 ( .o(net_9697), .ck(clk), .d(n3884) );
ms00f80  l0700 ( .o(net_9700), .ck(clk), .d(n3889) );
ms00f80  l0701 ( .o(_net_9363), .ck(clk), .d(n3894) );
ms00f80  l0702 ( .o(_net_190), .ck(clk), .d(n3899) );
ms00f80  l0703 ( .o(net_9747), .ck(clk), .d(n3904) );
ms00f80  l0704 ( .o(net_9840), .ck(clk), .d(n3909) );
ms00f80  l0705 ( .o(_net_10269), .ck(clk), .d(n3914) );
ms00f80  l0706 ( .o(net_9280), .ck(clk), .d(n3919) );
ms00f80  l0707 ( .o(net_245), .ck(clk), .d(n3923) );
ms00f80  l0708 ( .o(_net_10458), .ck(clk), .d(n3928) );
ms00f80  l0709 ( .o(net_289), .ck(clk), .d(n3933) );
ms00f80  l0710 ( .o(net_194), .ck(clk), .d(n3937) );
ms00f80  l0711 ( .o(_net_9161), .ck(clk), .d(n3942) );
ms00f80  l0712 ( .o(net_137), .ck(clk), .d(n3947) );
ms00f80  l0713 ( .o(net_10498), .ck(clk), .d(n3952) );
ms00f80  l0714 ( .o(net_9264), .ck(clk), .d(n3957) );
ms00f80  l0715 ( .o(net_9119), .ck(clk), .d(n3962) );
ms00f80  l0716 ( .o(_net_9187), .ck(clk), .d(n3967) );
ms00f80  l0717 ( .o(_net_10114), .ck(clk), .d(n3972) );
ms00f80  l0718 ( .o(x784), .ck(clk), .d(n3976) );
ms00f80  l0719 ( .o(_net_9356), .ck(clk), .d(n3980) );
ms00f80  l0720 ( .o(net_9973), .ck(clk), .d(n3985) );
ms00f80  l0721 ( .o(net_9288), .ck(clk), .d(n3990) );
ms00f80  l0722 ( .o(_net_9643), .ck(clk), .d(n3994) );
ms00f80  l0723 ( .o(_net_10151), .ck(clk), .d(n3999) );
ms00f80  l0724 ( .o(net_9760), .ck(clk), .d(n4004) );
ms00f80  l0725 ( .o(net_10133), .ck(clk), .d(n4009) );
ms00f80  l0726 ( .o(_net_10143), .ck(clk), .d(n4014) );
ms00f80  l0727 ( .o(net_9906), .ck(clk), .d(n4019) );
ms00f80  l0728 ( .o(_net_10109), .ck(clk), .d(n4024) );
ms00f80  l0729 ( .o(_net_10426), .ck(clk), .d(n4029) );
ms00f80  l0730 ( .o(_net_254), .ck(clk), .d(n4034) );
ms00f80  l0731 ( .o(net_9813), .ck(clk), .d(n4039) );
ms00f80  l0732 ( .o(net_9873), .ck(clk), .d(n4044) );
ms00f80  l0733 ( .o(_net_10334), .ck(clk), .d(n4049) );
ms00f80  l0734 ( .o(_net_10249), .ck(clk), .d(n4054) );
ms00f80  l0735 ( .o(net_223), .ck(clk), .d(n4059) );
ms00f80  l0736 ( .o(net_9270), .ck(clk), .d(n4064) );
ms00f80  l0737 ( .o(_net_10441), .ck(clk), .d(n4069) );
ms00f80  l0738 ( .o(net_10404), .ck(clk), .d(n4074) );
ms00f80  l0739 ( .o(net_9807), .ck(clk), .d(n4079) );
ms00f80  l0740 ( .o(net_9283), .ck(clk), .d(n4084) );
ms00f80  l0741 ( .o(_net_9557), .ck(clk), .d(n4088) );
ms00f80  l0742 ( .o(_net_10316), .ck(clk), .d(n4093) );
ms00f80  l0743 ( .o(net_9594), .ck(clk), .d(n4098) );
ms00f80  l0744 ( .o(net_9852), .ck(clk), .d(n4103) );
ms00f80  l0745 ( .o(net_9453), .ck(clk), .d(n4108) );
ms00f80  l0746 ( .o(_net_9250), .ck(clk), .d(n4112) );
ms00f80  l0747 ( .o(x1215), .ck(clk), .d(n4116) );
ms00f80  l0748 ( .o(net_9340), .ck(clk), .d(n4120) );
ms00f80  l0749 ( .o(net_9737), .ck(clk), .d(n4124) );
ms00f80  l0750 ( .o(_net_10480), .ck(clk), .d(n4129) );
ms00f80  l0751 ( .o(x454), .ck(clk), .d(n4133) );
ms00f80  l0752 ( .o(net_9718), .ck(clk), .d(n4137) );
ms00f80  l0753 ( .o(_net_9402), .ck(clk), .d(n4142) );
ms00f80  l0754 ( .o(net_10297), .ck(clk), .d(n4147) );
ms00f80  l0755 ( .o(net_9252), .ck(clk), .d(n4151) );
ms00f80  l0756 ( .o(net_9903), .ck(clk), .d(n4156) );
ms00f80  l0757 ( .o(net_114), .ck(clk), .d(n4161) );
ms00f80  l0758 ( .o(_net_9832), .ck(clk), .d(n4165) );
ms00f80  l0759 ( .o(_net_10250), .ck(clk), .d(n4170) );
ms00f80  l0760 ( .o(net_9841), .ck(clk), .d(n4175) );
ms00f80  l0761 ( .o(_net_121), .ck(clk), .d(n4180) );
ms00f80  l0762 ( .o(net_10067), .ck(clk), .d(n4185) );
ms00f80  l0763 ( .o(_net_8840), .ck(clk), .d(n4190) );
ms00f80  l0764 ( .o(net_9758), .ck(clk), .d(n4195) );
ms00f80  l0765 ( .o(_net_10346), .ck(clk), .d(n4200) );
ms00f80  l0766 ( .o(_net_10464), .ck(clk), .d(n4205) );
ms00f80  l0767 ( .o(_net_9232), .ck(clk), .d(n4210) );
ms00f80  l0768 ( .o(_net_10138), .ck(clk), .d(n4215) );
ms00f80  l0769 ( .o(_net_166), .ck(clk), .d(n4220) );
ms00f80  l0770 ( .o(_net_161), .ck(clk), .d(n4225) );
ms00f80  l0771 ( .o(net_10183), .ck(clk), .d(n4230) );
ms00f80  l0772 ( .o(_net_10146), .ck(clk), .d(n4235) );
ms00f80  l0773 ( .o(net_9529), .ck(clk), .d(n4240) );
ms00f80  l0774 ( .o(net_9892), .ck(clk), .d(n4245) );
ms00f80  l0775 ( .o(_net_10529), .ck(clk), .d(n4250) );
ms00f80  l0776 ( .o(net_301), .ck(clk), .d(n4255) );
ms00f80  l0777 ( .o(_net_9312), .ck(clk), .d(n4259) );
ms00f80  l0778 ( .o(_net_9602), .ck(clk), .d(n4264) );
ms00f80  l0779 ( .o(_net_10358), .ck(clk), .d(n4269) );
ms00f80  l0780 ( .o(net_113), .ck(clk), .d(n4274) );
ms00f80  l0781 ( .o(net_10408), .ck(clk), .d(n4279) );
ms00f80  l0782 ( .o(net_9269), .ck(clk), .d(n4283) );
ms00f80  l0783 ( .o(net_9657), .ck(clk), .d(n4288) );
ms00f80  l0784 ( .o(net_9631), .ck(clk), .d(n4293) );
ms00f80  l0785 ( .o(net_9149), .ck(clk), .d(n4298) );
ms00f80  l0786 ( .o(net_9776), .ck(clk), .d(n4303) );
ms00f80  l0787 ( .o(net_10023), .ck(clk), .d(n4308) );
ms00f80  l0788 ( .o(net_9357), .ck(clk), .d(n4312) );
ms00f80  l0789 ( .o(net_252), .ck(clk), .d(n4316) );
ms00f80  l0790 ( .o(net_9664), .ck(clk), .d(n4321) );
ms00f80  l0791 ( .o(net_10079), .ck(clk), .d(n4326) );
ms00f80  l0792 ( .o(_net_9296), .ck(clk), .d(n4331) );
ms00f80  l0793 ( .o(net_9872), .ck(clk), .d(n4336) );
ms00f80  l0794 ( .o(_net_9409), .ck(clk), .d(n4341) );
ms00f80  l0795 ( .o(_net_10255), .ck(clk), .d(n4346) );
ms00f80  l0796 ( .o(net_9260), .ck(clk), .d(n4351) );
ms00f80  l0797 ( .o(net_9759), .ck(clk), .d(n4355) );
ms00f80  l0798 ( .o(net_9584), .ck(clk), .d(n4360) );
ms00f80  l0799 ( .o(net_9465), .ck(clk), .d(n4364) );
ms00f80  l0800 ( .o(x1298), .ck(clk), .d(n4368) );
ms00f80  l0801 ( .o(_net_9949), .ck(clk), .d(n4372) );
ms00f80  l0802 ( .o(net_9964), .ck(clk), .d(n4377) );
ms00f80  l0803 ( .o(net_9597), .ck(clk), .d(n4382) );
ms00f80  l0804 ( .o(net_9534), .ck(clk), .d(n4387) );
ms00f80  l0805 ( .o(_net_9941), .ck(clk), .d(n4392) );
ms00f80  l0806 ( .o(net_10019), .ck(clk), .d(n4397) );
ms00f80  l0807 ( .o(x871), .ck(clk), .d(n4401) );
ms00f80  l0808 ( .o(_net_10339), .ck(clk), .d(n4405) );
ms00f80  l0809 ( .o(net_9128), .ck(clk), .d(n4410) );
ms00f80  l0810 ( .o(_net_10475), .ck(clk), .d(n4415) );
ms00f80  l0811 ( .o(_net_233), .ck(clk), .d(n4420) );
ms00f80  l0812 ( .o(_net_9243), .ck(clk), .d(n4425) );
ms00f80  l0813 ( .o(x1343), .ck(clk), .d(n4430) );
ms00f80  l0814 ( .o(net_9780), .ck(clk), .d(n4434) );
ms00f80  l0815 ( .o(_net_167), .ck(clk), .d(n4439) );
ms00f80  l0816 ( .o(net_9889), .ck(clk), .d(n4444) );
ms00f80  l0817 ( .o(net_9682), .ck(clk), .d(n4449) );
ms00f80  l0818 ( .o(net_9670), .ck(clk), .d(n4454) );
ms00f80  l0819 ( .o(_net_10153), .ck(clk), .d(n4459) );
ms00f80  l0820 ( .o(net_10514), .ck(clk), .d(n4463) );
ms00f80  l0821 ( .o(_net_9411), .ck(clk), .d(n4468) );
ms00f80  l0822 ( .o(net_203), .ck(clk), .d(n4473) );
ms00f80  l0823 ( .o(net_9497), .ck(clk), .d(n4477) );
ms00f80  l0824 ( .o(net_10283), .ck(clk), .d(n4482) );
ms00f80  l0825 ( .o(_net_9541), .ck(clk), .d(n4487) );
ms00f80  l0826 ( .o(_net_9196), .ck(clk), .d(n4491) );
ms00f80  l0827 ( .o(net_10300), .ck(clk), .d(n4496) );
ms00f80  l0828 ( .o(net_10281), .ck(clk), .d(n4501) );
ms00f80  l0829 ( .o(net_9919), .ck(clk), .d(n4506) );
ms00f80  l0830 ( .o(_net_171), .ck(clk), .d(n4511) );
ms00f80  l0831 ( .o(_net_10341), .ck(clk), .d(n4516) );
ms00f80  l0832 ( .o(x1074), .ck(clk), .d(n4521) );
ms00f80  l0833 ( .o(net_9918), .ck(clk), .d(n4525) );
ms00f80  l0834 ( .o(net_10010), .ck(clk), .d(n4530) );
ms00f80  l0835 ( .o(net_306), .ck(clk), .d(n4535) );
ms00f80  l0836 ( .o(_net_8830), .ck(clk), .d(n4539) );
ms00f80  l0837 ( .o(_net_154), .ck(clk), .d(n4544) );
ms00f80  l0838 ( .o(net_9308), .ck(clk), .d(n4549) );
ms00f80  l0839 ( .o(net_9809), .ck(clk), .d(n4554) );
ms00f80  l0840 ( .o(net_9685), .ck(clk), .d(n4559) );
ms00f80  l0841 ( .o(_net_10340), .ck(clk), .d(n4564) );
ms00f80  l0842 ( .o(net_9698), .ck(clk), .d(n4569) );
ms00f80  l0843 ( .o(net_9124), .ck(clk), .d(n4574) );
ms00f80  l0844 ( .o(_net_9572), .ck(clk), .d(n4579) );
ms00f80  l0845 ( .o(net_10523), .ck(clk), .d(n4584) );
ms00f80  l0846 ( .o(_net_10196), .ck(clk), .d(n4589) );
ms00f80  l0847 ( .o(_net_120), .ck(clk), .d(n4594) );
ms00f80  l0848 ( .o(net_9568), .ck(clk), .d(n4598) );
ms00f80  l0849 ( .o(net_10082), .ck(clk), .d(n4603) );
ms00f80  l0850 ( .o(_net_9839), .ck(clk), .d(n4608) );
ms00f80  l0851 ( .o(_net_10279), .ck(clk), .d(n4613) );
ms00f80  l0852 ( .o(net_9847), .ck(clk), .d(n4618) );
ms00f80  l0853 ( .o(_net_10202), .ck(clk), .d(n4623) );
ms00f80  l0854 ( .o(net_9262), .ck(clk), .d(n4627) );
ms00f80  l0855 ( .o(_net_9645), .ck(clk), .d(n4632) );
ms00f80  l0856 ( .o(net_10398), .ck(clk), .d(n4637) );
ms00f80  l0857 ( .o(_net_9611), .ck(clk), .d(n4642) );
ms00f80  l0858 ( .o(net_292), .ck(clk), .d(n4647) );
ms00f80  l0859 ( .o(x1282), .ck(clk), .d(n4650) );
ms00f80  l0860 ( .o(net_9907), .ck(clk), .d(n4654) );
ms00f80  l0861 ( .o(net_209), .ck(clk), .d(n4659) );
ms00f80  l0862 ( .o(_net_10430), .ck(clk), .d(n4664) );
ms00f80  l0863 ( .o(_net_9547), .ck(clk), .d(n4668) );
ms00f80  l0864 ( .o(net_9703), .ck(clk), .d(n4673) );
ms00f80  l0865 ( .o(net_10274), .ck(clk), .d(n4678) );
ms00f80  l0866 ( .o(net_10199), .ck(clk), .d(n4682) );
ms00f80  l0867 ( .o(_net_9406), .ck(clk), .d(n4687) );
ms00f80  l0868 ( .o(net_295), .ck(clk), .d(n4692) );
ms00f80  l0869 ( .o(net_9210), .ck(clk), .d(n4696) );
ms00f80  l0870 ( .o(net_9559), .ck(clk), .d(n4700) );
ms00f80  l0871 ( .o(net_10015), .ck(clk), .d(n4705) );
ms00f80  l0872 ( .o(_net_178), .ck(clk), .d(n4710) );
ms00f80  l0873 ( .o(x962), .ck(clk), .d(n4715) );
ms00f80  l0874 ( .o(net_10185), .ck(clk), .d(n4719) );
ms00f80  l0875 ( .o(_net_8847), .ck(clk), .d(n4724) );
ms00f80  l0876 ( .o(net_10051), .ck(clk), .d(n4729) );
ms00f80  l0877 ( .o(_net_10148), .ck(clk), .d(n4734) );
ms00f80  l0878 ( .o(net_144), .ck(clk), .d(n4739) );
ms00f80  l0879 ( .o(net_9513), .ck(clk), .d(n4744) );
ms00f80  l0880 ( .o(_net_9215), .ck(clk), .d(n4749) );
ms00f80  l0881 ( .o(net_9613), .ck(clk), .d(n4754) );
ms00f80  l0882 ( .o(net_9755), .ck(clk), .d(n4759) );
ms00f80  l0883 ( .o(net_9696), .ck(clk), .d(n4764) );
ms00f80  l0884 ( .o(_net_10265), .ck(clk), .d(n4769) );
ms00f80  l0885 ( .o(net_9617), .ck(clk), .d(n4774) );
ms00f80  l0886 ( .o(net_9896), .ck(clk), .d(n4779) );
ms00f80  l0887 ( .o(net_297), .ck(clk), .d(n4784) );
ms00f80  l0888 ( .o(net_9882), .ck(clk), .d(n4788) );
ms00f80  l0889 ( .o(net_9659), .ck(clk), .d(n4793) );
ms00f80  l0890 ( .o(net_9216), .ck(clk), .d(n4797) );
ms00f80  l0891 ( .o(net_9858), .ck(clk), .d(n4802) );
ms00f80  l0892 ( .o(_net_151), .ck(clk), .d(n4807) );
ms00f80  l0893 ( .o(_net_10120), .ck(clk), .d(n4812) );
ms00f80  l0894 ( .o(net_9920), .ck(clk), .d(n4817) );
ms00f80  l0895 ( .o(net_9787), .ck(clk), .d(n4822) );
ms00f80  l0896 ( .o(net_10052), .ck(clk), .d(n4827) );
ms00f80  l0897 ( .o(net_9936), .ck(clk), .d(n4832) );
ms00f80  l0898 ( .o(net_9975), .ck(clk), .d(n4837) );
ms00f80  l0899 ( .o(x1248), .ck(clk), .d(n4842) );
ms00f80  l0900 ( .o(net_10003), .ck(clk), .d(n4846) );
ms00f80  l0901 ( .o(_net_10117), .ck(clk), .d(n4851) );
ms00f80  l0902 ( .o(_net_9415), .ck(clk), .d(n4856) );
ms00f80  l0903 ( .o(net_236), .ck(clk), .d(n4861) );
ms00f80  l0904 ( .o(net_9683), .ck(clk), .d(n4866) );
ms00f80  l0905 ( .o(_net_9519), .ck(clk), .d(n4871) );
ms00f80  l0906 ( .o(net_95), .ck(clk), .d(n4875) );
ms00f80  l0907 ( .o(net_10286), .ck(clk), .d(n4879) );
ms00f80  l0908 ( .o(net_10080), .ck(clk), .d(n4884) );
ms00f80  l0909 ( .o(_net_9566), .ck(clk), .d(n4889) );
ms00f80  l0910 ( .o(_net_10383), .ck(clk), .d(n4894) );
ms00f80  l0911 ( .o(_net_174), .ck(clk), .d(n4899) );
ms00f80  l0912 ( .o(net_10517), .ck(clk), .d(n4904) );
ms00f80  l0913 ( .o(net_216), .ck(clk), .d(n4908) );
ms00f80  l0914 ( .o(_net_10112), .ck(clk), .d(n4913) );
ms00f80  l0915 ( .o(net_9836), .ck(clk), .d(n4918) );
ms00f80  l0916 ( .o(_net_9169), .ck(clk), .d(n4923) );
ms00f80  l0917 ( .o(_net_9040), .ck(clk), .d(n4927) );
ms00f80  l0918 ( .o(_net_9311), .ck(clk), .d(n4932) );
ms00f80  l0919 ( .o(x526), .ck(clk), .d(n4937) );
ms00f80  l0920 ( .o(net_10022), .ck(clk), .d(n4941) );
ms00f80  l0921 ( .o(_net_10515), .ck(clk), .d(n4946) );
ms00f80  l0922 ( .o(net_9668), .ck(clk), .d(n4951) );
ms00f80  l0923 ( .o(net_9968), .ck(clk), .d(n4956) );
ms00f80  l0924 ( .o(_net_10355), .ck(clk), .d(n4961) );
ms00f80  l0925 ( .o(net_9197), .ck(clk), .d(n4966) );
ms00f80  l0926 ( .o(_net_10145), .ck(clk), .d(n4971) );
ms00f80  l0927 ( .o(net_308), .ck(clk), .d(n4976) );
ms00f80  l0928 ( .o(net_9884), .ck(clk), .d(n4980) );
ms00f80  l0929 ( .o(_net_10204), .ck(clk), .d(n4985) );
ms00f80  l0930 ( .o(_net_10418), .ck(clk), .d(n4990) );
ms00f80  l0931 ( .o(net_9436), .ck(clk), .d(n4995) );
ms00f80  l0932 ( .o(_net_9646), .ck(clk), .d(n5000) );
ms00f80  l0933 ( .o(_net_9309), .ck(clk), .d(n5005) );
ms00f80  l0934 ( .o(net_10397), .ck(clk), .d(n5010) );
ms00f80  l0935 ( .o(_net_10173), .ck(clk), .d(n5015) );
ms00f80  l0936 ( .o(_net_10324), .ck(clk), .d(n5020) );
ms00f80  l0937 ( .o(_net_9395), .ck(clk), .d(n5025) );
ms00f80  l0938 ( .o(net_9795), .ck(clk), .d(n5030) );
ms00f80  l0939 ( .o(net_10541), .ck(clk), .d(n5035) );
ms00f80  l0940 ( .o(net_10527), .ck(clk), .d(n5038) );
ms00f80  l0941 ( .o(_net_10471), .ck(clk), .d(n5043) );
ms00f80  l0942 ( .o(_net_10428), .ck(clk), .d(n5048) );
ms00f80  l0943 ( .o(net_9233), .ck(clk), .d(n5052) );
ms00f80  l0944 ( .o(_net_10172), .ck(clk), .d(n5057) );
ms00f80  l0945 ( .o(net_229), .ck(clk), .d(n5062) );
ms00f80  l0946 ( .o(net_10089), .ck(clk), .d(n5067) );
ms00f80  l0947 ( .o(net_9993), .ck(clk), .d(n5072) );
ms00f80  l0948 ( .o(net_9765), .ck(clk), .d(n5077) );
ms00f80  l0949 ( .o(net_9279), .ck(clk), .d(n5082) );
ms00f80  l0950 ( .o(net_9304), .ck(clk), .d(n5087) );
ms00f80  l0951 ( .o(net_9727), .ck(clk), .d(n5091) );
ms00f80  l0952 ( .o(_net_10056), .ck(clk), .d(n5096) );
ms00f80  l0953 ( .o(net_9282), .ck(clk), .d(n5101) );
ms00f80  l0954 ( .o(net_9762), .ck(clk), .d(n5105) );
ms00f80  l0955 ( .o(net_9692), .ck(clk), .d(n5110) );
ms00f80  l0956 ( .o(_net_9326), .ck(clk), .d(n5115) );
ms00f80  l0957 ( .o(_net_10062), .ck(clk), .d(n5120) );
ms00f80  l0958 ( .o(_net_9929), .ck(clk), .d(n5125) );
ms00f80  l0959 ( .o(_net_10465), .ck(clk), .d(n5130) );
ms00f80  l0960 ( .o(net_9890), .ck(clk), .d(n5135) );
ms00f80  l0961 ( .o(x1231), .ck(clk), .d(n5139) );
ms00f80  l0962 ( .o(_net_9391), .ck(clk), .d(n5143) );
ms00f80  l0963 ( .o(_net_9258), .ck(clk), .d(n5147) );
ms00f80  l0964 ( .o(net_9701), .ck(clk), .d(n5152) );
ms00f80  l0965 ( .o(net_9445), .ck(clk), .d(n5157) );
ms00f80  l0966 ( .o(net_9327), .ck(clk), .d(n5161) );
ms00f80  l0967 ( .o(net_9464), .ck(clk), .d(n5165) );
ms00f80  l0968 ( .o(_net_9740), .ck(clk), .d(n5169) );
ms00f80  l0969 ( .o(net_9676), .ck(clk), .d(n5174) );
ms00f80  l0970 ( .o(_net_10161), .ck(clk), .d(n5179) );
ms00f80  l0971 ( .o(_net_10469), .ck(clk), .d(n5184) );
ms00f80  l0972 ( .o(_net_10337), .ck(clk), .d(n5189) );
ms00f80  l0973 ( .o(net_304), .ck(clk), .d(n5194) );
ms00f80  l0974 ( .o(net_9822), .ck(clk), .d(n5198) );
ms00f80  l0975 ( .o(net_111), .ck(clk), .d(n5203) );
ms00f80  l0976 ( .o(_net_10235), .ck(clk), .d(n5208) );
ms00f80  l0977 ( .o(net_9498), .ck(clk), .d(n5212) );
ms00f80  l0978 ( .o(_net_9416), .ck(clk), .d(n5217) );
ms00f80  l0979 ( .o(net_9121), .ck(clk), .d(n5222) );
ms00f80  l0980 ( .o(net_207), .ck(clk), .d(n5227) );
ms00f80  l0981 ( .o(net_9271), .ck(clk), .d(n5232) );
ms00f80  l0982 ( .o(net_9914), .ck(clk), .d(n5237) );
ms00f80  l0983 ( .o(_net_10460), .ck(clk), .d(n5242) );
ms00f80  l0984 ( .o(net_9714), .ck(clk), .d(n5247) );
ms00f80  l0985 ( .o(net_150), .ck(clk), .d(n5252) );
ms00f80  l0986 ( .o(net_9768), .ck(clk), .d(n5257) );
ms00f80  l0987 ( .o(net_298), .ck(clk), .d(n5262) );
ms00f80  l0988 ( .o(x1313), .ck(clk), .d(n5266) );
ms00f80  l0989 ( .o(_net_162), .ck(clk), .d(n5270) );
ms00f80  l0990 ( .o(net_9369), .ck(clk), .d(n5275) );
ms00f80  l0991 ( .o(x1187), .ck(clk), .d(n5279) );
ms00f80  l0992 ( .o(_net_9628), .ck(clk), .d(n5283) );
ms00f80  l0993 ( .o(_net_277), .ck(clk), .d(n5288) );
ms00f80  l0994 ( .o(_net_276), .ck(clk), .d(n5293) );
ms00f80  l0995 ( .o(net_96), .ck(clk), .d(n5297) );
ms00f80  l0996 ( .o(_net_132), .ck(clk), .d(n5302) );
ms00f80  l0997 ( .o(_net_10197), .ck(clk), .d(n5306) );
ms00f80  l0998 ( .o(_net_175), .ck(clk), .d(n5311) );
ms00f80  l0999 ( .o(_net_10124), .ck(clk), .d(n5316) );
ms00f80  l1000 ( .o(_net_10164), .ck(clk), .d(n5321) );
ms00f80  l1001 ( .o(_net_10245), .ck(clk), .d(n5326) );
ms00f80  l1002 ( .o(_net_9399), .ck(clk), .d(n5331) );
ms00f80  l1003 ( .o(_net_9209), .ck(clk), .d(n5336) );
ms00f80  l1004 ( .o(_net_10463), .ck(clk), .d(n5341) );
ms00f80  l1005 ( .o(net_9837), .ck(clk), .d(n5346) );
ms00f80  l1006 ( .o(x1142), .ck(clk), .d(n5351) );
ms00f80  l1007 ( .o(net_10063), .ck(clk), .d(n5355) );
ms00f80  l1008 ( .o(net_9666), .ck(clk), .d(n5360) );
ms00f80  l1009 ( .o(net_204), .ck(clk), .d(n5365) );
ms00f80  l1010 ( .o(net_9358), .ck(clk), .d(n5370) );
ms00f80  l1011 ( .o(net_9339), .ck(clk), .d(n5375) );
ms00f80  l1012 ( .o(net_9793), .ck(clk), .d(n5379) );
ms00f80  l1013 ( .o(_net_182), .ck(clk), .d(n5384) );
ms00f80  l1014 ( .o(net_9857), .ck(clk), .d(n5389) );
ms00f80  l1015 ( .o(_net_10141), .ck(clk), .d(n5394) );
ms00f80  l1016 ( .o(_net_126), .ck(clk), .d(n5399) );
ms00f80  l1017 ( .o(net_10537), .ck(clk), .d(n5403) );
ms00f80  l1018 ( .o(net_9285), .ck(clk), .d(n5408) );
ms00f80  l1019 ( .o(_net_10119), .ck(clk), .d(n5412) );
ms00f80  l1020 ( .o(net_9365), .ck(clk), .d(n5417) );
ms00f80  l1021 ( .o(net_8820), .ck(clk), .d(n5422) );
ms00f80  l1022 ( .o(_net_10159), .ck(clk), .d(n5427) );
ms00f80  l1023 ( .o(net_9549), .ck(clk), .d(n5431) );
ms00f80  l1024 ( .o(_net_10360), .ck(clk), .d(n5436) );
ms00f80  l1025 ( .o(_net_9588), .ck(clk), .d(n5441) );
ms00f80  l1026 ( .o(_net_8869), .ck(clk), .d(n5445) );
ms00f80  l1027 ( .o(_net_9268), .ck(clk), .d(n5449) );
ms00f80  l1028 ( .o(net_9705), .ck(clk), .d(n5454) );
ms00f80  l1029 ( .o(_net_10370), .ck(clk), .d(n5459) );
ms00f80  l1030 ( .o(_net_9407), .ck(clk), .d(n5464) );
ms00f80  l1031 ( .o(net_9136), .ck(clk), .d(n5469) );
ms00f80  l1032 ( .o(net_9448), .ck(clk), .d(n5473) );
ms00f80  l1033 ( .o(net_9329), .ck(clk), .d(n5477) );
ms00f80  l1034 ( .o(net_10402), .ck(clk), .d(n5481) );
ms00f80  l1035 ( .o(_net_10338), .ck(clk), .d(n5486) );
ms00f80  l1036 ( .o(_net_272), .ck(clk), .d(n5491) );
ms00f80  l1037 ( .o(_net_9558), .ck(clk), .d(n5495) );
ms00f80  l1038 ( .o(_net_9728), .ck(clk), .d(n5500) );
ms00f80  l1039 ( .o(net_94), .ck(clk), .d(n5504) );
ms00f80  l1040 ( .o(net_9508), .ck(clk), .d(n5508) );
ms00f80  l1041 ( .o(net_9989), .ck(clk), .d(n5513) );
ms00f80  l1042 ( .o(net_9569), .ck(clk), .d(n5518) );
ms00f80  l1043 ( .o(_net_10305), .ck(clk), .d(n5523) );
ms00f80  l1044 ( .o(net_9289), .ck(clk), .d(n5528) );
ms00f80  l1045 ( .o(net_9150), .ck(clk), .d(n5533) );
ms00f80  l1046 ( .o(_net_10263), .ck(clk), .d(n5537) );
ms00f80  l1047 ( .o(_net_10438), .ck(clk), .d(n5542) );
ms00f80  l1048 ( .o(_net_9393), .ck(clk), .d(n5547) );
ms00f80  l1049 ( .o(_net_180), .ck(clk), .d(n5552) );
ms00f80  l1050 ( .o(net_9854), .ck(clk), .d(n5557) );
ms00f80  l1051 ( .o(_net_193), .ck(clk), .d(n5562) );
ms00f80  l1052 ( .o(_net_10354), .ck(clk), .d(n5567) );
ms00f80  l1053 ( .o(net_9615), .ck(clk), .d(n5572) );
ms00f80  l1054 ( .o(_net_9627), .ck(clk), .d(n5577) );
ms00f80  l1055 ( .o(net_288), .ck(clk), .d(n5582) );
ms00f80  l1056 ( .o(net_9153), .ck(clk), .d(n5585) );
ms00f80  l1057 ( .o(net_9485), .ck(clk), .d(n5589) );
ms00f80  l1058 ( .o(net_290), .ck(clk), .d(n5594) );
ms00f80  l1059 ( .o(net_98), .ck(clk), .d(n5597) );
ms00f80  l1060 ( .o(net_9449), .ck(clk), .d(n5601) );
ms00f80  l1061 ( .o(net_9278), .ck(clk), .d(n5605) );
ms00f80  l1062 ( .o(_net_10425), .ck(clk), .d(n5610) );
ms00f80  l1063 ( .o(net_9499), .ck(clk), .d(n5614) );
ms00f80  l1064 ( .o(net_10014), .ck(clk), .d(n5619) );
ms00f80  l1065 ( .o(net_9876), .ck(clk), .d(n5624) );
ms00f80  l1066 ( .o(net_9469), .ck(clk), .d(n5629) );
ms00f80  l1067 ( .o(_net_9661), .ck(clk), .d(n5633) );
ms00f80  l1068 ( .o(net_9335), .ck(clk), .d(n5638) );
ms00f80  l1069 ( .o(_net_156), .ck(clk), .d(n5642) );
ms00f80  l1070 ( .o(net_10018), .ck(clk), .d(n5647) );
ms00f80  l1071 ( .o(net_9257), .ck(clk), .d(n5651) );
ms00f80  l1072 ( .o(_net_9173), .ck(clk), .d(n5656) );
ms00f80  l1073 ( .o(_net_234), .ck(clk), .d(n5661) );
ms00f80  l1074 ( .o(_net_10212), .ck(clk), .d(n5666) );
ms00f80  l1075 ( .o(net_9713), .ck(clk), .d(n5671) );
ms00f80  l1076 ( .o(_net_9166), .ck(clk), .d(n5676) );
ms00f80  l1077 ( .o(net_294), .ck(clk), .d(n5681) );
ms00f80  l1078 ( .o(net_10066), .ck(clk), .d(n5685) );
ms00f80  l1079 ( .o(_net_8955), .ck(clk), .d(n5690) );
ms00f80  l1080 ( .o(_net_9928), .ck(clk), .d(n5695) );
ms00f80  l1081 ( .o(_net_9374), .ck(clk), .d(n5700) );
ms00f80  l1082 ( .o(net_10237), .ck(clk), .d(n5705) );
ms00f80  l1083 ( .o(net_10379), .ck(clk), .d(n5710) );
ms00f80  l1084 ( .o(net_9480), .ck(clk), .d(n5714) );
ms00f80  l1085 ( .o(net_242), .ck(clk), .d(n5719) );
ms00f80  l1086 ( .o(_net_10377), .ck(clk), .d(n5724) );
ms00f80  l1087 ( .o(net_10386), .ck(clk), .d(n5729) );
ms00f80  l1088 ( .o(net_102), .ck(clk), .d(n5734) );
ms00f80  l1089 ( .o(_net_9537), .ck(clk), .d(n5739) );
ms00f80  l1090 ( .o(x1010), .ck(clk), .d(n5744) );
ms00f80  l1091 ( .o(_net_10166), .ck(clk), .d(n5748) );
ms00f80  l1092 ( .o(_net_9324), .ck(clk), .d(n5753) );
ms00f80  l1093 ( .o(_net_10320), .ck(clk), .d(n5758) );
ms00f80  l1094 ( .o(net_9764), .ck(clk), .d(n5763) );
ms00f80  l1095 ( .o(_net_10042), .ck(clk), .d(n5768) );
ms00f80  l1096 ( .o(_net_10419), .ck(clk), .d(n5773) );
ms00f80  l1097 ( .o(net_240), .ck(clk), .d(n5777) );
ms00f80  l1098 ( .o(net_10285), .ck(clk), .d(n5782) );
ms00f80  l1099 ( .o(net_9966), .ck(clk), .d(n5787) );
ms00f80  l1100 ( .o(_net_9638), .ck(clk), .d(n5792) );
ms00f80  l1101 ( .o(net_9877), .ck(clk), .d(n5797) );
ms00f80  l1102 ( .o(net_10046), .ck(clk), .d(n5802) );
ms00f80  l1103 ( .o(_net_9355), .ck(clk), .d(n5807) );
ms00f80  l1104 ( .o(net_9336), .ck(clk), .d(n5812) );
ms00f80  l1105 ( .o(_net_9503), .ck(clk), .d(n5815) );
ms00f80  l1106 ( .o(_net_10277), .ck(clk), .d(n5820) );
ms00f80  l1107 ( .o(_net_10350), .ck(clk), .d(n5825) );
ms00f80  l1108 ( .o(_net_9520), .ck(clk), .d(n5830) );
ms00f80  l1109 ( .o(net_9144), .ck(clk), .d(n5835) );
ms00f80  l1110 ( .o(net_9868), .ck(clk), .d(n5839) );
ms00f80  l1111 ( .o(_net_9345), .ck(clk), .d(n5844) );
ms00f80  l1112 ( .o(_net_9398), .ck(clk), .d(n5849) );
ms00f80  l1113 ( .o(net_9542), .ck(clk), .d(n5853) );
ms00f80  l1114 ( .o(net_9432), .ck(clk), .d(n5858) );
ms00f80  l1115 ( .o(net_9887), .ck(clk), .d(n5863) );
ms00f80  l1116 ( .o(_net_9178), .ck(clk), .d(n5868) );
ms00f80  l1117 ( .o(_net_10130), .ck(clk), .d(n5873) );
ms00f80  l1118 ( .o(_net_10221), .ck(clk), .d(n5878) );
ms00f80  l1119 ( .o(net_9707), .ck(clk), .d(n5883) );
ms00f80  l1120 ( .o(_net_10412), .ck(clk), .d(n5888) );
ms00f80  l1121 ( .o(net_9980), .ck(clk), .d(n5893) );
ms00f80  l1122 ( .o(_net_10097), .ck(clk), .d(n5898) );
ms00f80  l1123 ( .o(_net_9957), .ck(clk), .d(n5903) );
ms00f80  l1124 ( .o(_net_10102), .ck(clk), .d(n5908) );
ms00f80  l1125 ( .o(_net_10261), .ck(clk), .d(n5913) );
ms00f80  l1126 ( .o(net_9152), .ck(clk), .d(n5917) );
ms00f80  l1127 ( .o(net_10083), .ck(clk), .d(n5921) );
ms00f80  l1128 ( .o(net_9783), .ck(clk), .d(n5926) );
ms00f80  l1129 ( .o(_net_10260), .ck(clk), .d(n5931) );
ms00f80  l1130 ( .o(net_9507), .ck(clk), .d(n5935) );
ms00f80  l1131 ( .o(net_9506), .ck(clk), .d(n5939) );
ms00f80  l1132 ( .o(net_230), .ck(clk), .d(n5944) );
ms00f80  l1133 ( .o(net_9711), .ck(clk), .d(n5949) );
ms00f80  l1134 ( .o(net_9726), .ck(clk), .d(n5954) );
ms00f80  l1135 ( .o(_net_10481), .ck(clk), .d(n5959) );
ms00f80  l1136 ( .o(net_9806), .ck(clk), .d(n5964) );
ms00f80  l1137 ( .o(net_241), .ck(clk), .d(n5969) );
ms00f80  l1138 ( .o(x1192), .ck(clk), .d(n5974) );
ms00f80  l1139 ( .o(net_212), .ck(clk), .d(n5978) );
ms00f80  l1140 ( .o(net_9571), .ck(clk), .d(n5983) );
ms00f80  l1141 ( .o(net_10509), .ck(clk), .d(n5988) );
ms00f80  l1142 ( .o(net_9772), .ck(clk), .d(n5993) );
ms00f80  l1143 ( .o(net_9334), .ck(clk), .d(n5998) );
ms00f80  l1144 ( .o(net_10516), .ck(clk), .d(n6001) );
ms00f80  l1145 ( .o(net_279), .ck(clk), .d(n6005) );
ms00f80  l1146 ( .o(x1402), .ck(clk), .d(n6009) );
ms00f80  l1147 ( .o(net_8837), .ck(clk), .d(n6013) );
ms00f80  l1148 ( .o(_net_10140), .ck(clk), .d(n6018) );
ms00f80  l1149 ( .o(_net_10057), .ck(clk), .d(n6023) );
ms00f80  l1150 ( .o(net_9689), .ck(clk), .d(n6028) );
ms00f80  l1151 ( .o(net_9163), .ck(clk), .d(n6033) );
ms00f80  l1152 ( .o(_net_9203), .ck(clk), .d(n6037) );
ms00f80  l1153 ( .o(_net_10462), .ck(clk), .d(n6042) );
ms00f80  l1154 ( .o(net_9526), .ck(clk), .d(n6047) );
ms00f80  l1155 ( .o(_net_201), .ck(clk), .d(n6052) );
ms00f80  l1156 ( .o(_net_160), .ck(clk), .d(n6057) );
ms00f80  l1157 ( .o(_net_9833), .ck(clk), .d(n6062) );
ms00f80  l1158 ( .o(net_9251), .ck(clk), .d(n6067) );
ms00f80  l1159 ( .o(_net_176), .ck(clk), .d(n6072) );
ms00f80  l1160 ( .o(net_10510), .ck(clk), .d(n6077) );
ms00f80  l1161 ( .o(net_9866), .ck(clk), .d(n6082) );
ms00f80  l1162 ( .o(net_147), .ck(clk), .d(n6087) );
ms00f80  l1163 ( .o(net_300), .ck(clk), .d(n6091) );
ms00f80  l1164 ( .o(net_9462), .ck(clk), .d(n6095) );
ms00f80  l1165 ( .o(net_9467), .ck(clk), .d(n6099) );
ms00f80  l1166 ( .o(_net_9546), .ck(clk), .d(n6102) );
ms00f80  l1167 ( .o(net_9131), .ck(clk), .d(n6107) );
ms00f80  l1168 ( .o(net_9721), .ck(clk), .d(n6111) );
ms00f80  l1169 ( .o(_net_10424), .ck(clk), .d(n6116) );
ms00f80  l1170 ( .o(net_10342), .ck(clk), .d(n6121) );
ms00f80  l1171 ( .o(net_9784), .ck(clk), .d(n6126) );
ms00f80  l1172 ( .o(net_9425), .ck(clk), .d(n6131) );
ms00f80  l1173 ( .o(net_9200), .ck(clk), .d(n6136) );
ms00f80  l1174 ( .o(net_10345), .ck(clk), .d(n6141) );
ms00f80  l1175 ( .o(net_238), .ck(clk), .d(n6145) );
ms00f80  l1176 ( .o(_net_10456), .ck(clk), .d(n6150) );
ms00f80  l1177 ( .o(_net_10367), .ck(clk), .d(n6155) );
ms00f80  l1178 ( .o(net_139), .ck(clk), .d(n6160) );
ms00f80  l1179 ( .o(_net_189), .ck(clk), .d(n6164) );
ms00f80  l1180 ( .o(net_9287), .ck(clk), .d(n6169) );
ms00f80  l1181 ( .o(_net_9752), .ck(clk), .d(n6173) );
ms00f80  l1182 ( .o(net_10525), .ck(clk), .d(n6177) );
ms00f80  l1183 ( .o(net_9261), .ck(clk), .d(n6181) );
ms00f80  l1184 ( .o(_net_10444), .ck(clk), .d(n6186) );
ms00f80  l1185 ( .o(_net_9734), .ck(clk), .d(n6191) );
ms00f80  l1186 ( .o(net_10191), .ck(clk), .d(n6196) );
ms00f80  l1187 ( .o(net_10134), .ck(clk), .d(n6201) );
ms00f80  l1188 ( .o(_net_9934), .ck(clk), .d(n6206) );
ms00f80  l1189 ( .o(net_9977), .ck(clk), .d(n6211) );
ms00f80  l1190 ( .o(_net_9299), .ck(clk), .d(n6216) );
ms00f80  l1191 ( .o(_net_10037), .ck(clk), .d(n6221) );
ms00f80  l1192 ( .o(net_9838), .ck(clk), .d(n6226) );
ms00f80  l1193 ( .o(net_10170), .ck(clk), .d(n6231) );
ms00f80  l1194 ( .o(net_10524), .ck(clk), .d(n6235) );
ms00f80  l1195 ( .o(net_283), .ck(clk), .d(n6240) );
ms00f80  l1196 ( .o(_net_10457), .ck(clk), .d(n6244) );
ms00f80  l1197 ( .o(net_10044), .ck(clk), .d(n6249) );
ms00f80  l1198 ( .o(x1274), .ck(clk), .d(n6254) );
ms00f80  l1199 ( .o(net_9699), .ck(clk), .d(n6258) );
ms00f80  l1200 ( .o(_net_10416), .ck(clk), .d(n6263) );
ms00f80  l1201 ( .o(_net_10026), .ck(clk), .d(n6268) );
ms00f80  l1202 ( .o(net_93), .ck(clk), .d(n6272) );
ms00f80  l1203 ( .o(_net_10321), .ck(clk), .d(n6277) );
ms00f80  l1204 ( .o(_net_9944), .ck(clk), .d(n6282) );
ms00f80  l1205 ( .o(_net_10442), .ck(clk), .d(n6287) );
ms00f80  l1206 ( .o(net_9991), .ck(clk), .d(n6292) );
ms00f80  l1207 ( .o(net_9535), .ck(clk), .d(n6297) );
ms00f80  l1208 ( .o(net_9442), .ck(clk), .d(n6302) );
ms00f80  l1209 ( .o(_net_9239), .ck(clk), .d(n6306) );
ms00f80  l1210 ( .o(_net_9422), .ck(clk), .d(n6311) );
ms00f80  l1211 ( .o(net_9716), .ck(clk), .d(n6316) );
ms00f80  l1212 ( .o(net_10403), .ck(clk), .d(n6321) );
ms00f80  l1213 ( .o(net_9766), .ck(clk), .d(n6326) );
ms00f80  l1214 ( .o(_net_10325), .ck(clk), .d(n6331) );
ms00f80  l1215 ( .o(net_8827), .ck(clk), .d(n6336) );
ms00f80  l1216 ( .o(net_9674), .ck(clk), .d(n6341) );
ms00f80  l1217 ( .o(net_9757), .ck(clk), .d(n6346) );
ms00f80  l1218 ( .o(_net_9413), .ck(clk), .d(n6351) );
ms00f80  l1219 ( .o(net_9138), .ck(clk), .d(n6356) );
ms00f80  l1220 ( .o(net_9331), .ck(clk), .d(n6360) );
ms00f80  l1221 ( .o(_net_261), .ck(clk), .d(n6364) );
ms00f80  l1222 ( .o(net_9306), .ck(clk), .d(n6369) );
ms00f80  l1223 ( .o(net_9946), .ck(clk), .d(n6373) );
ms00f80  l1224 ( .o(net_9935), .ck(clk), .d(n6378) );
ms00f80  l1225 ( .o(_net_10259), .ck(clk), .d(n6383) );
ms00f80  l1226 ( .o(_net_9423), .ck(clk), .d(n6388) );
ms00f80  l1227 ( .o(net_9126), .ck(clk), .d(n6393) );
ms00f80  l1228 ( .o(net_9596), .ck(clk), .d(n6397) );
ms00f80  l1229 ( .o(_net_9556), .ck(clk), .d(n6401) );
ms00f80  l1230 ( .o(net_9982), .ck(clk), .d(n6406) );
ms00f80  l1231 ( .o(_net_10207), .ck(clk), .d(n6411) );
ms00f80  l1232 ( .o(_net_10427), .ck(clk), .d(n6416) );
ms00f80  l1233 ( .o(_net_10128), .ck(clk), .d(n6421) );
ms00f80  l1234 ( .o(_net_9293), .ck(clk), .d(n6426) );
ms00f80  l1235 ( .o(net_9923), .ck(clk), .d(n6431) );
ms00f80  l1236 ( .o(_net_9168), .ck(clk), .d(n6436) );
ms00f80  l1237 ( .o(_net_10310), .ck(clk), .d(n6441) );
ms00f80  l1238 ( .o(net_10405), .ck(clk), .d(n6446) );
ms00f80  l1239 ( .o(net_148), .ck(clk), .d(n6451) );
ms00f80  l1240 ( .o(_net_9401), .ck(clk), .d(n6456) );
ms00f80  l1241 ( .o(net_9470), .ck(clk), .d(n6460) );
ms00f80  l1242 ( .o(net_9477), .ck(clk), .d(n6464) );
ms00f80  l1243 ( .o(net_10495), .ck(clk), .d(n6469) );
ms00f80  l1244 ( .o(net_9349), .ck(clk), .d(n6474) );
ms00f80  l1245 ( .o(net_10000), .ck(clk), .d(n6479) );
ms00f80  l1246 ( .o(_net_10230), .ck(clk), .d(n6484) );
ms00f80  l1247 ( .o(_net_10215), .ck(clk), .d(n6489) );
ms00f80  l1248 ( .o(net_9490), .ck(clk), .d(n6493) );
ms00f80  l1249 ( .o(net_9803), .ck(clk), .d(n6498) );
ms00f80  l1250 ( .o(_net_10111), .ck(clk), .d(n6503) );
ms00f80  l1251 ( .o(net_9478), .ck(clk), .d(n6507) );
ms00f80  l1252 ( .o(net_9531), .ck(clk), .d(n6512) );
ms00f80  l1253 ( .o(_net_9403), .ck(clk), .d(n6517) );
ms00f80  l1254 ( .o(x637), .ck(clk), .d(n6522) );
ms00f80  l1255 ( .o(net_9742), .ck(clk), .d(n6526) );
ms00f80  l1256 ( .o(_net_10329), .ck(clk), .d(n6531) );
ms00f80  l1257 ( .o(_net_123), .ck(clk), .d(n6536) );
ms00f80  l1258 ( .o(_net_9235), .ck(clk), .d(n6541) );
ms00f80  l1259 ( .o(_net_118), .ck(clk), .d(n6546) );
ms00f80  l1260 ( .o(net_9969), .ck(clk), .d(n6551) );
ms00f80  l1261 ( .o(_net_9376), .ck(clk), .d(n6556) );
ms00f80  l1262 ( .o(net_10069), .ck(clk), .d(n6561) );
ms00f80  l1263 ( .o(_net_9207), .ck(clk), .d(n6566) );
ms00f80  l1264 ( .o(net_9148), .ck(clk), .d(n6571) );
ms00f80  l1265 ( .o(net_9777), .ck(clk), .d(n6575) );
ms00f80  l1266 ( .o(net_9491), .ck(clk), .d(n6579) );
ms00f80  l1267 ( .o(net_247), .ck(clk), .d(n6584) );
ms00f80  l1268 ( .o(net_9812), .ck(clk), .d(n6589) );
ms00f80  l1269 ( .o(_net_9515), .ck(clk), .d(n6594) );
ms00f80  l1270 ( .o(net_9864), .ck(clk), .d(n6599) );
ms00f80  l1271 ( .o(_net_271), .ck(clk), .d(n6604) );
ms00f80  l1272 ( .o(net_9753), .ck(clk), .d(n6609) );
ms00f80  l1273 ( .o(net_9223), .ck(clk), .d(n6614) );
ms00f80  l1274 ( .o(net_220), .ck(clk), .d(n6619) );
ms00f80  l1275 ( .o(_net_10474), .ck(clk), .d(n6624) );
ms00f80  l1276 ( .o(_net_188), .ck(clk), .d(n6629) );
ms00f80  l1277 ( .o(net_9648), .ck(clk), .d(n6634) );
ms00f80  l1278 ( .o(net_10289), .ck(clk), .d(n6639) );
ms00f80  l1279 ( .o(_net_10171), .ck(clk), .d(n6644) );
ms00f80  l1280 ( .o(_net_10030), .ck(clk), .d(n6649) );
ms00f80  l1281 ( .o(_net_159), .ck(clk), .d(n6654) );
ms00f80  l1282 ( .o(net_9899), .ck(clk), .d(n6659) );
ms00f80  l1283 ( .o(net_8816), .ck(clk), .d(n6664) );
ms00f80  l1284 ( .o(_net_10095), .ck(clk), .d(n6669) );
ms00f80  l1285 ( .o(_net_10155), .ck(clk), .d(n6674) );
ms00f80  l1286 ( .o(_net_10364), .ck(clk), .d(n6679) );
ms00f80  l1287 ( .o(net_9725), .ck(clk), .d(n6684) );
ms00f80  l1288 ( .o(net_226), .ck(clk), .d(n6689) );
ms00f80  l1289 ( .o(net_10344), .ck(clk), .d(n6694) );
ms00f80  l1290 ( .o(_net_8819), .ck(clk), .d(n6699) );
ms00f80  l1291 ( .o(net_9348), .ck(clk), .d(n6704) );
ms00f80  l1292 ( .o(_net_9427), .ck(clk), .d(n6709) );
ms00f80  l1293 ( .o(net_9475), .ck(clk), .d(n6713) );
ms00f80  l1294 ( .o(_net_9567), .ck(clk), .d(n6718) );
ms00f80  l1295 ( .o(_net_10244), .ck(clk), .d(n6723) );
ms00f80  l1296 ( .o(_net_9958), .ck(clk), .d(n6728) );
ms00f80  l1297 ( .o(net_146), .ck(clk), .d(n6733) );
ms00f80  l1298 ( .o(net_10491), .ck(clk), .d(n6738) );
ms00f80  l1299 ( .o(net_9754), .ck(clk), .d(n6743) );
ms00f80  l1300 ( .o(net_9622), .ck(clk), .d(n6748) );
ms00f80  l1301 ( .o(net_9667), .ck(clk), .d(n6753) );
ms00f80  l1302 ( .o(_net_10121), .ck(clk), .d(n6758) );
ms00f80  l1303 ( .o(_net_9564), .ck(clk), .d(n6763) );
ms00f80  l1304 ( .o(net_9781), .ck(clk), .d(n6768) );
ms00f80  l1305 ( .o(net_9179), .ck(clk), .d(n6773) );
ms00f80  l1306 ( .o(_net_179), .ck(clk), .d(n6778) );
ms00f80  l1307 ( .o(x1153), .ck(clk), .d(n6782) );
ms00f80  l1308 ( .o(net_10399), .ck(clk), .d(n6786) );
ms00f80  l1309 ( .o(net_9791), .ck(clk), .d(n6791) );
ms00f80  l1310 ( .o(net_9690), .ck(clk), .d(n6796) );
ms00f80  l1311 ( .o(net_9865), .ck(clk), .d(n6801) );
ms00f80  l1312 ( .o(net_9771), .ck(clk), .d(n6806) );
ms00f80  l1313 ( .o(_net_173), .ck(clk), .d(n6811) );
ms00f80  l1314 ( .o(net_260), .ck(clk), .d(n6816) );
ms00f80  l1315 ( .o(net_10085), .ck(clk), .d(n6821) );
ms00f80  l1316 ( .o(_net_9845), .ck(clk), .d(n6826) );
ms00f80  l1317 ( .o(net_9796), .ck(clk), .d(n6831) );
ms00f80  l1318 ( .o(net_9624), .ck(clk), .d(n6836) );
ms00f80  l1319 ( .o(net_142), .ck(clk), .d(n6841) );
ms00f80  l1320 ( .o(_net_10165), .ck(clk), .d(n6846) );
ms00f80  l1321 ( .o(net_9675), .ck(clk), .d(n6851) );
ms00f80  l1322 ( .o(_net_9297), .ck(clk), .d(n6856) );
ms00f80  l1323 ( .o(_net_9851), .ck(clk), .d(n6861) );
ms00f80  l1324 ( .o(net_9170), .ck(clk), .d(n6865) );
ms00f80  l1325 ( .o(_net_10157), .ck(clk), .d(n6870) );
ms00f80  l1326 ( .o(_net_10234), .ck(clk), .d(n6875) );
ms00f80  l1327 ( .o(_net_10246), .ck(clk), .d(n6880) );
ms00f80  l1328 ( .o(net_9574), .ck(clk), .d(n6885) );
ms00f80  l1329 ( .o(net_10004), .ck(clk), .d(n6890) );
ms00f80  l1330 ( .o(_net_9176), .ck(clk), .d(n6895) );
ms00f80  l1331 ( .o(_net_10439), .ck(clk), .d(n6900) );
ms00f80  l1332 ( .o(_net_10032), .ck(clk), .d(n6905) );
ms00f80  l1333 ( .o(x1384), .ck(clk), .d(n6910) );
ms00f80  l1334 ( .o(net_9663), .ck(clk), .d(n6914) );
ms00f80  l1335 ( .o(_net_9384), .ck(clk), .d(n6919) );
ms00f80  l1336 ( .o(_net_10118), .ck(clk), .d(n6924) );
ms00f80  l1337 ( .o(_net_10381), .ck(clk), .d(n6929) );
ms00f80  l1338 ( .o(net_10401), .ck(clk), .d(n6934) );
ms00f80  l1339 ( .o(net_10485), .ck(clk), .d(n6939) );
ms00f80  l1340 ( .o(_net_9266), .ck(clk), .d(n6944) );
ms00f80  l1341 ( .o(_net_9532), .ck(clk), .d(n6949) );
ms00f80  l1342 ( .o(net_9145), .ck(clk), .d(n6954) );
ms00f80  l1343 ( .o(net_251), .ck(clk), .d(n6958) );
ms00f80  l1344 ( .o(net_257), .ck(clk), .d(n6962) );
ms00f80  l1345 ( .o(net_9472), .ck(clk), .d(n6966) );
ms00f80  l1346 ( .o(_net_10241), .ck(clk), .d(n6971) );
ms00f80  l1347 ( .o(_net_10208), .ck(clk), .d(n6976) );
ms00f80  l1348 ( .o(x987), .ck(clk), .d(n6981) );
ms00f80  l1349 ( .o(net_9440), .ck(clk), .d(n6985) );
ms00f80  l1350 ( .o(net_9820), .ck(clk), .d(n6989) );
ms00f80  l1351 ( .o(net_9254), .ck(clk), .d(n6993) );
ms00f80  l1352 ( .o(net_10070), .ck(clk), .d(n6998) );
ms00f80  l1353 ( .o(net_9623), .ck(clk), .d(n7003) );
ms00f80  l1354 ( .o(net_91), .ck(clk), .d(n7007) );
ms00f80  l1355 ( .o(_net_10152), .ck(clk), .d(n7012) );
ms00f80  l1356 ( .o(_net_10330), .ck(clk), .d(n7017) );
ms00f80  l1357 ( .o(_net_10407), .ck(clk), .d(n7021) );
ms00f80  l1358 ( .o(net_10288), .ck(clk), .d(n7026) );
ms00f80  l1359 ( .o(net_9156), .ck(clk), .d(n7030) );
ms00f80  l1360 ( .o(net_10075), .ck(clk), .d(n7034) );
ms00f80  l1361 ( .o(net_10287), .ck(clk), .d(n7039) );
ms00f80  l1362 ( .o(net_9455), .ck(clk), .d(n7044) );
ms00f80  l1363 ( .o(net_9798), .ck(clk), .d(n7048) );
ms00f80  l1364 ( .o(_net_255), .ck(clk), .d(n7053) );
ms00f80  l1365 ( .o(net_9651), .ck(clk), .d(n7058) );
ms00f80  l1366 ( .o(net_9276), .ck(clk), .d(n7063) );
ms00f80  l1367 ( .o(_net_9295), .ck(clk), .d(n7068) );
ms00f80  l1368 ( .o(_net_9189), .ck(clk), .d(n7073) );
ms00f80  l1369 ( .o(net_291), .ck(clk), .d(n7078) );
ms00f80  l1370 ( .o(net_10293), .ck(clk), .d(n7082) );
ms00f80  l1371 ( .o(net_248), .ck(clk), .d(n7086) );
ms00f80  l1372 ( .o(net_9756), .ck(clk), .d(n7091) );
ms00f80  l1373 ( .o(_net_9551), .ck(clk), .d(n7095) );
ms00f80  l1374 ( .o(net_9458), .ck(clk), .d(n7100) );
ms00f80  l1375 ( .o(_net_9412), .ck(clk), .d(n7104) );
ms00f80  l1376 ( .o(_net_10094), .ck(clk), .d(n7108) );
ms00f80  l1377 ( .o(net_9778), .ck(clk), .d(n7113) );
ms00f80  l1378 ( .o(_net_10041), .ck(clk), .d(n7118) );
ms00f80  l1379 ( .o(net_9789), .ck(clk), .d(n7123) );
ms00f80  l1380 ( .o(_net_10433), .ck(clk), .d(n7128) );
ms00f80  l1381 ( .o(net_10074), .ck(clk), .d(n7133) );
ms00f80  l1382 ( .o(_net_10099), .ck(clk), .d(n7138) );
ms00f80  l1383 ( .o(_net_10486), .ck(clk), .d(n7143) );
ms00f80  l1384 ( .o(net_9704), .ck(clk), .d(n7148) );
ms00f80  l1385 ( .o(net_9805), .ck(clk), .d(n7153) );
ms00f80  l1386 ( .o(net_9598), .ck(clk), .d(n7158) );
ms00f80  l1387 ( .o(net_9431), .ck(clk), .d(n7163) );
ms00f80  l1388 ( .o(_net_10160), .ck(clk), .d(n7168) );
ms00f80  l1389 ( .o(net_9141), .ck(clk), .d(n7173) );
ms00f80  l1390 ( .o(net_9222), .ck(clk), .d(n7177) );
ms00f80  l1391 ( .o(net_10389), .ck(clk), .d(n7182) );
ms00f80  l1392 ( .o(_net_10043), .ck(clk), .d(n7187) );
ms00f80  l1393 ( .o(net_9702), .ck(clk), .d(n7192) );
ms00f80  l1394 ( .o(_net_280), .ck(clk), .d(n7197) );
ms00f80  l1395 ( .o(_net_10200), .ck(clk), .d(n7202) );
ms00f80  l1396 ( .o(net_10304), .ck(clk), .d(n7206) );
ms00f80  l1397 ( .o(_net_9658), .ck(clk), .d(n7211) );
ms00f80  l1398 ( .o(net_9855), .ck(clk), .d(n7216) );
ms00f80  l1399 ( .o(_net_9397), .ck(clk), .d(n7221) );
ms00f80  l1400 ( .o(_net_9352), .ck(clk), .d(n7226) );
ms00f80  l1401 ( .o(net_9125), .ck(clk), .d(n7231) );
ms00f80  l1402 ( .o(net_10035), .ck(clk), .d(n7235) );
ms00f80  l1403 ( .o(net_9671), .ck(clk), .d(n7240) );
ms00f80  l1404 ( .o(net_9874), .ck(clk), .d(n7245) );
ms00f80  l1405 ( .o(net_10036), .ck(clk), .d(n7250) );
ms00f80  l1406 ( .o(net_10184), .ck(clk), .d(n7255) );
ms00f80  l1407 ( .o(_net_8834), .ck(clk), .d(n7260) );
ms00f80  l1408 ( .o(_net_9290), .ck(clk), .d(n7265) );
ms00f80  l1409 ( .o(_net_10236), .ck(clk), .d(n7270) );
ms00f80  l1410 ( .o(net_9693), .ck(clk), .d(n7275) );
ms00f80  l1411 ( .o(net_9681), .ck(clk), .d(n7280) );
ms00f80  l1412 ( .o(net_9763), .ck(clk), .d(n7285) );
ms00f80  l1413 ( .o(net_10504), .ck(clk), .d(n7290) );
ms00f80  l1414 ( .o(_net_198), .ck(clk), .d(n7295) );
ms00f80  l1415 ( .o(net_9225), .ck(clk), .d(n7300) );
ms00f80  l1416 ( .o(x1262), .ck(clk), .d(n7304) );
ms00f80  l1417 ( .o(net_10198), .ck(clk), .d(n7308) );
ms00f80  l1418 ( .o(_net_9516), .ck(clk), .d(n7312) );
ms00f80  l1419 ( .o(net_9307), .ck(clk), .d(n7317) );
ms00f80  l1420 ( .o(_net_10437), .ck(clk), .d(n7321) );
ms00f80  l1421 ( .o(net_10492), .ck(clk), .d(n7326) );
ms00f80  l1422 ( .o(net_9971), .ck(clk), .d(n7331) );
ms00f80  l1423 ( .o(net_10282), .ck(clk), .d(n7336) );
ms00f80  l1424 ( .o(_net_170), .ck(clk), .d(n7341) );
ms00f80  l1425 ( .o(net_10396), .ck(clk), .d(n7346) );
ms00f80  l1426 ( .o(_net_10168), .ck(clk), .d(n7351) );
ms00f80  l1427 ( .o(net_195), .ck(clk), .d(n7355) );
ms00f80  l1428 ( .o(net_9976), .ck(clk), .d(n7360) );
ms00f80  l1429 ( .o(_net_9636), .ck(clk), .d(n7365) );
ms00f80  l1430 ( .o(net_227), .ck(clk), .d(n7370) );
ms00f80  l1431 ( .o(net_134), .ck(clk), .d(n7375) );
ms00f80  l1432 ( .o(net_9219), .ck(clk), .d(n7379) );
ms00f80  l1433 ( .o(net_10188), .ck(clk), .d(n7384) );
ms00f80  l1434 ( .o(net_9961), .ck(clk), .d(n7389) );
ms00f80  l1435 ( .o(net_9593), .ck(clk), .d(n7394) );
ms00f80  l1436 ( .o(_net_9555), .ck(clk), .d(n7398) );
ms00f80  l1437 ( .o(net_9985), .ck(clk), .d(n7403) );
ms00f80  l1438 ( .o(net_186), .ck(clk), .d(n7408) );
ms00f80  l1439 ( .o(_net_10314), .ck(clk), .d(n7413) );
ms00f80  l1440 ( .o(net_9632), .ck(clk), .d(n7418) );
ms00f80  l1441 ( .o(_net_10445), .ck(clk), .d(n7423) );
ms00f80  l1442 ( .o(net_143), .ck(clk), .d(n7428) );
ms00f80  l1443 ( .o(_net_8821), .ck(clk), .d(n7432) );
ms00f80  l1444 ( .o(net_9501), .ck(clk), .d(n7436) );
ms00f80  l1445 ( .o(net_9231), .ck(clk), .d(n7441) );
ms00f80  l1446 ( .o(_net_9378), .ck(clk), .d(n7446) );
ms00f80  l1447 ( .o(net_138), .ck(clk), .d(n7451) );
ms00f80  l1448 ( .o(_net_10228), .ck(clk), .d(n7455) );
ms00f80  l1449 ( .o(net_9987), .ck(clk), .d(n7460) );
ms00f80  l1450 ( .o(_net_199), .ck(clk), .d(n7465) );
ms00f80  l1451 ( .o(_net_9429), .ck(clk), .d(n7470) );
ms00f80  l1452 ( .o(_net_9301), .ck(clk), .d(n7475) );
ms00f80  l1453 ( .o(net_9450), .ck(clk), .d(n7480) );
ms00f80  l1454 ( .o(_net_9746), .ck(clk), .d(n7484) );
ms00f80  l1455 ( .o(net_9198), .ck(clk), .d(n7489) );
ms00f80  l1456 ( .o(net_9861), .ck(clk), .d(n7494) );
ms00f80  l1457 ( .o(_net_10272), .ck(clk), .d(n7499) );
ms00f80  l1458 ( .o(net_10076), .ck(clk), .d(n7504) );
ms00f80  l1459 ( .o(net_10400), .ck(clk), .d(n7509) );
ms00f80  l1460 ( .o(net_10071), .ck(clk), .d(n7514) );
ms00f80  l1461 ( .o(net_9997), .ck(clk), .d(n7519) );
ms00f80  l1462 ( .o(net_10500), .ck(clk), .d(n7524) );
ms00f80  l1463 ( .o(net_10391), .ck(clk), .d(n7529) );
ms00f80  l1464 ( .o(net_9586), .ck(clk), .d(n7534) );
ms00f80  l1465 ( .o(net_9494), .ck(clk), .d(n7538) );
ms00f80  l1466 ( .o(_net_10459), .ck(clk), .d(n7543) );
ms00f80  l1467 ( .o(x769), .ck(clk), .d(n7548) );
ms00f80  l1468 ( .o(_net_9214), .ck(clk), .d(n7552) );
ms00f80  l1469 ( .o(net_10280), .ck(clk), .d(n7557) );
ms00f80  l1470 ( .o(x1029), .ck(clk), .d(n7562) );
ms00f80  l1471 ( .o(_net_10267), .ck(clk), .d(n7566) );
ms00f80  l1472 ( .o(_net_10306), .ck(clk), .d(n7571) );
ms00f80  l1473 ( .o(net_9482), .ck(clk), .d(n7575) );
ms00f80  l1474 ( .o(net_243), .ck(clk), .d(n7580) );
ms00f80  l1475 ( .o(net_9885), .ck(clk), .d(n7585) );
ms00f80  l1476 ( .o(net_10385), .ck(clk), .d(n7590) );
ms00f80  l1477 ( .o(net_110), .ck(clk), .d(n7595) );
ms00f80  l1478 ( .o(net_9739), .ck(clk), .d(n7600) );
ms00f80  l1479 ( .o(net_105), .ck(clk), .d(n7605) );
ms00f80  l1480 ( .o(net_9719), .ck(clk), .d(n7609) );
ms00f80  l1481 ( .o(x1104), .ck(clk), .d(n7613) );
ms00f80  l1482 ( .o(net_9444), .ck(clk), .d(n7617) );
ms00f80  l1483 ( .o(_net_9418), .ck(clk), .d(n7621) );
ms00f80  l1484 ( .o(_net_10332), .ck(clk), .d(n7626) );
ms00f80  l1485 ( .o(net_222), .ck(clk), .d(n7631) );
ms00f80  l1486 ( .o(net_9910), .ck(clk), .d(n7636) );
ms00f80  l1487 ( .o(net_9476), .ck(clk), .d(n7640) );
ms00f80  l1488 ( .o(net_10505), .ck(clk), .d(n7645) );
ms00f80  l1489 ( .o(_net_10472), .ck(clk), .d(n7650) );
ms00f80  l1490 ( .o(_net_9926), .ck(clk), .d(n7655) );
ms00f80  l1491 ( .o(_net_9204), .ck(clk), .d(n7660) );
ms00f80  l1492 ( .o(_net_9842), .ck(clk), .d(n7665) );
ms00f80  l1493 ( .o(net_205), .ck(clk), .d(n7670) );
ms00f80  l1494 ( .o(net_10532), .ck(clk), .d(n7675) );
ms00f80  l1495 ( .o(net_9709), .ck(clk), .d(n7680) );
ms00f80  l1496 ( .o(net_9953), .ck(clk), .d(n7685) );
ms00f80  l1497 ( .o(_net_177), .ck(clk), .d(n7690) );
ms00f80  l1498 ( .o(_net_9635), .ck(clk), .d(n7695) );
ms00f80  l1499 ( .o(_net_10268), .ck(clk), .d(n7700) );
ms00f80  l1500 ( .o(net_237), .ck(clk), .d(n7704) );
ms00f80  l1501 ( .o(net_9310), .ck(clk), .d(n7709) );
ms00f80  l1502 ( .o(_net_9353), .ck(clk), .d(n7714) );
ms00f80  l1503 ( .o(_net_9389), .ck(clk), .d(n7719) );
ms00f80  l1504 ( .o(net_10238), .ck(clk), .d(n7724) );
ms00f80  l1505 ( .o(_net_10106), .ck(clk), .d(n7729) );
ms00f80  l1506 ( .o(net_286), .ck(clk), .d(n7734) );
ms00f80  l1507 ( .o(_net_10466), .ck(clk), .d(n7738) );
ms00f80  l1508 ( .o(_net_9733), .ck(clk), .d(n7743) );
ms00f80  l1509 ( .o(net_10449), .ck(clk), .d(n7748) );
ms00f80  l1510 ( .o(_net_9240), .ck(clk), .d(n7753) );
ms00f80  l1511 ( .o(_net_10454), .ck(clk), .d(n7758) );
ms00f80  l1512 ( .o(net_8832), .ck(clk), .d(n7763) );
ms00f80  l1513 ( .o(_net_10422), .ck(clk), .d(n7768) );
ms00f80  l1514 ( .o(_net_10455), .ck(clk), .d(n7773) );
ms00f80  l1515 ( .o(net_9368), .ck(clk), .d(n7778) );
ms00f80  l1516 ( .o(_net_9548), .ck(clk), .d(n7782) );
ms00f80  l1517 ( .o(_net_10327), .ck(clk), .d(n7787) );
ms00f80  l1518 ( .o(net_9120), .ck(clk), .d(n7792) );
ms00f80  l1519 ( .o(_net_9373), .ck(clk), .d(n7796) );
ms00f80  l1520 ( .o(net_10298), .ck(clk), .d(n7801) );
ms00f80  l1521 ( .o(_net_200), .ck(clk), .d(n7806) );
ms00f80  l1522 ( .o(_net_10254), .ck(clk), .d(n7811) );
ms00f80  l1523 ( .o(_net_9730), .ck(clk), .d(n7816) );
ms00f80  l1524 ( .o(_net_10423), .ck(clk), .d(n7821) );
ms00f80  l1525 ( .o(net_9974), .ck(clk), .d(n7826) );
ms00f80  l1526 ( .o(x1329), .ck(clk), .d(n7830) );
ms00f80  l1527 ( .o(_net_10415), .ck(clk), .d(n7834) );
ms00f80  l1528 ( .o(net_9123), .ck(clk), .d(n7839) );
ms00f80  l1529 ( .o(net_9706), .ck(clk), .d(n7843) );
ms00f80  l1530 ( .o(_net_9388), .ck(clk), .d(n7848) );
ms00f80  l1531 ( .o(net_9147), .ck(clk), .d(n7853) );
ms00f80  l1532 ( .o(_net_9321), .ck(clk), .d(n7857) );
ms00f80  l1533 ( .o(net_303), .ck(clk), .d(n7862) );
ms00f80  l1534 ( .o(_net_9603), .ck(clk), .d(n7866) );
ms00f80  l1535 ( .o(_net_9732), .ck(clk), .d(n7871) );
ms00f80  l1536 ( .o(_net_10476), .ck(clk), .d(n7876) );
ms00f80  l1537 ( .o(net_9817), .ck(clk), .d(n7881) );
ms00f80  l1538 ( .o(net_9259), .ck(clk), .d(n7885) );
ms00f80  l1539 ( .o(net_115), .ck(clk), .d(n7889) );
ms00f80  l1540 ( .o(net_235), .ck(clk), .d(n7893) );
ms00f80  l1541 ( .o(net_9925), .ck(clk), .d(n7898) );
ms00f80  l1542 ( .o(net_9361), .ck(clk), .d(n7902) );
ms00f80  l1543 ( .o(_net_9381), .ck(clk), .d(n7906) );
ms00f80  l1544 ( .o(net_9875), .ck(clk), .d(n7911) );
ms00f80  l1545 ( .o(_net_9421), .ck(clk), .d(n7916) );
ms00f80  l1546 ( .o(_net_10055), .ck(clk), .d(n7921) );
ms00f80  l1547 ( .o(net_10522), .ck(clk), .d(n7925) );
ms00f80  l1548 ( .o(net_10024), .ck(clk), .d(n7930) );
ms00f80  l1549 ( .o(net_10012), .ck(clk), .d(n7935) );
ms00f80  l1550 ( .o(net_10078), .ck(clk), .d(n7940) );
ms00f80  l1551 ( .o(_net_8826), .ck(clk), .d(n7945) );
ms00f80  l1552 ( .o(net_9129), .ck(clk), .d(n7950) );
ms00f80  l1553 ( .o(net_9457), .ck(clk), .d(n7954) );
ms00f80  l1554 ( .o(net_9509), .ck(clk), .d(n7957) );
ms00f80  l1555 ( .o(net_10169), .ck(clk), .d(n7962) );
ms00f80  l1556 ( .o(_net_10538), .ck(clk), .d(n7967) );
ms00f80  l1557 ( .o(_net_9428), .ck(clk), .d(n7972) );
ms00f80  l1558 ( .o(_net_10147), .ck(clk), .d(n7977) );
ms00f80  l1559 ( .o(net_9895), .ck(clk), .d(n7982) );
ms00f80  l1560 ( .o(net_9959), .ck(clk), .d(n7987) );
ms00f80  l1561 ( .o(net_10542), .ck(clk), .d(n7992) );
ms00f80  l1562 ( .o(_net_129), .ck(clk), .d(n7996) );
ms00f80  l1563 ( .o(_net_9521), .ck(clk), .d(n8001) );
ms00f80  l1564 ( .o(_net_164), .ck(clk), .d(n8006) );
ms00f80  l1565 ( .o(net_9539), .ck(clk), .d(n8011) );
ms00f80  l1566 ( .o(_net_10535), .ck(clk), .d(n8016) );
ms00f80  l1567 ( .o(_net_9609), .ck(clk), .d(n8021) );
ms00f80  l1568 ( .o(_net_232), .ck(clk), .d(n8026) );
ms00f80  l1569 ( .o(_net_10201), .ck(clk), .d(n8031) );
ms00f80  l1570 ( .o(net_10292), .ck(clk), .d(n8036) );
ms00f80  l1571 ( .o(_net_9843), .ck(clk), .d(n8041) );
ms00f80  l1572 ( .o(_net_9950), .ck(clk), .d(n8046) );
ms00f80  l1573 ( .o(_net_10322), .ck(clk), .d(n8051) );
ms00f80  l1574 ( .o(net_9263), .ck(clk), .d(n8055) );
ms00f80  l1575 ( .o(net_10177), .ck(clk), .d(n8059) );
ms00f80  l1576 ( .o(net_253), .ck(clk), .d(n8063) );
ms00f80  l1577 ( .o(net_9474), .ck(clk), .d(n8067) );
ms00f80  l1578 ( .o(net_9426), .ck(clk), .d(n8072) );
ms00f80  l1579 ( .o(net_10521), .ck(clk), .d(n8076) );
ms00f80  l1580 ( .o(net_9904), .ck(clk), .d(n8081) );
ms00f80  l1581 ( .o(_net_9291), .ck(clk), .d(n8086) );
ms00f80  l1582 ( .o(net_10013), .ck(clk), .d(n8091) );
ms00f80  l1583 ( .o(_net_9405), .ck(clk), .d(n8096) );
ms00f80  l1584 ( .o(net_9810), .ck(clk), .d(n8101) );
ms00f80  l1585 ( .o(_net_10131), .ck(clk), .d(n8106) );
ms00f80  l1586 ( .o(net_9779), .ck(clk), .d(n8111) );
ms00f80  l1587 ( .o(_net_9392), .ck(clk), .d(n8116) );
ms00f80  l1588 ( .o(net_9511), .ck(clk), .d(n8120) );
ms00f80  l1589 ( .o(net_9979), .ck(clk), .d(n8125) );
ms00f80  l1590 ( .o(_net_10105), .ck(clk), .d(n8130) );
ms00f80  l1591 ( .o(_net_9165), .ck(clk), .d(n8135) );
ms00f80  l1592 ( .o(_net_9316), .ck(clk), .d(n8140) );
ms00f80  l1593 ( .o(_net_10251), .ck(clk), .d(n8145) );
ms00f80  l1594 ( .o(_net_10301), .ck(clk), .d(n8150) );
ms00f80  l1595 ( .o(_net_9248), .ck(clk), .d(n8155) );
ms00f80  l1596 ( .o(net_9612), .ck(clk), .d(n8160) );
ms00f80  l1597 ( .o(_net_10421), .ck(clk), .d(n8165) );
ms00f80  l1598 ( .o(net_9853), .ck(clk), .d(n8170) );
ms00f80  l1599 ( .o(_net_10315), .ck(clk), .d(n8175) );
ms00f80  l1600 ( .o(net_10087), .ck(clk), .d(n8180) );
ms00f80  l1601 ( .o(net_9174), .ck(clk), .d(n8185) );
ms00f80  l1602 ( .o(net_9799), .ck(clk), .d(n8190) );
ms00f80  l1603 ( .o(net_9686), .ck(clk), .d(n8195) );
ms00f80  l1604 ( .o(_net_9408), .ck(clk), .d(n8200) );
ms00f80  l1605 ( .o(_net_9410), .ck(clk), .d(n8205) );
ms00f80  l1606 ( .o(net_10513), .ck(clk), .d(n8210) );
ms00f80  l1607 ( .o(net_10182), .ck(clk), .d(n8214) );
ms00f80  l1608 ( .o(net_9447), .ck(clk), .d(n8219) );
ms00f80  l1609 ( .o(_net_10142), .ck(clk), .d(n8223) );
ms00f80  l1610 ( .o(x1370), .ck(clk), .d(n8227) );
ms00f80  l1611 ( .o(net_9870), .ck(clk), .d(n8231) );
ms00f80  l1612 ( .o(_net_9550), .ck(clk), .d(n8235) );
ms00f80  l1613 ( .o(net_9909), .ck(clk), .d(n8240) );
ms00f80  l1614 ( .o(_net_9942), .ck(clk), .d(n8245) );
ms00f80  l1615 ( .o(_net_10049), .ck(clk), .d(n8250) );
ms00f80  l1616 ( .o(net_10186), .ck(clk), .d(n8255) );
ms00f80  l1617 ( .o(_net_10276), .ck(clk), .d(n8260) );
ms00f80  l1618 ( .o(x461), .ck(clk), .d(n8264) );
ms00f80  l1619 ( .o(_net_10270), .ck(clk), .d(n8268) );
ms00f80  l1620 ( .o(x1161), .ck(clk), .d(n8272) );
ms00f80  l1621 ( .o(net_10395), .ck(clk), .d(n8276) );
ms00f80  l1622 ( .o(net_10017), .ck(clk), .d(n8281) );
ms00f80  l1623 ( .o(net_9277), .ck(clk), .d(n8286) );
ms00f80  l1624 ( .o(_net_10213), .ck(clk), .d(n8291) );
ms00f80  l1625 ( .o(net_9999), .ck(clk), .d(n8296) );
ms00f80  l1626 ( .o(_net_133), .ck(clk), .d(n8301) );
ms00f80  l1627 ( .o(_net_10302), .ck(clk), .d(n8305) );
ms00f80  l1628 ( .o(net_10053), .ck(clk), .d(n8310) );
ms00f80  l1629 ( .o(_net_9211), .ck(clk), .d(n8315) );
ms00f80  l1630 ( .o(net_9770), .ck(clk), .d(n8320) );
ms00f80  l1631 ( .o(net_9863), .ck(clk), .d(n8325) );
ms00f80  l1632 ( .o(_net_9343), .ck(clk), .d(n8330) );
ms00f80  l1633 ( .o(net_10187), .ck(clk), .d(n8335) );
ms00f80  l1634 ( .o(net_10540), .ck(clk), .d(n8339) );
ms00f80  l1635 ( .o(net_10447), .ck(clk), .d(n8344) );
ms00f80  l1636 ( .o(net_9741), .ck(clk), .d(n8349) );
ms00f80  l1637 ( .o(net_112), .ck(clk), .d(n8354) );
ms00f80  l1638 ( .o(net_9720), .ck(clk), .d(n8358) );
ms00f80  l1639 ( .o(_net_10233), .ck(clk), .d(n8363) );
ms00f80  l1640 ( .o(net_293), .ck(clk), .d(n8368) );
ms00f80  l1641 ( .o(_net_10214), .ck(clk), .d(n8372) );
ms00f80  l1642 ( .o(net_9510), .ck(clk), .d(n8376) );
ms00f80  l1643 ( .o(net_9157), .ck(clk), .d(n8380) );
ms00f80  l1644 ( .o(net_9430), .ck(clk), .d(n8384) );
ms00f80  l1645 ( .o(net_219), .ck(clk), .d(n8389) );
ms00f80  l1646 ( .o(_net_10257), .ck(clk), .d(n8394) );
ms00f80  l1647 ( .o(_net_10278), .ck(clk), .d(n8399) );
ms00f80  l1648 ( .o(net_8835), .ck(clk), .d(n8404) );
ms00f80  l1649 ( .o(_net_9217), .ck(clk), .d(n8409) );
ms00f80  l1650 ( .o(net_224), .ck(clk), .d(n8414) );
ms00f80  l1651 ( .o(net_9797), .ck(clk), .d(n8419) );
ms00f80  l1652 ( .o(_net_153), .ck(clk), .d(n8424) );
ms00f80  l1653 ( .o(net_9599), .ck(clk), .d(n8429) );
ms00f80  l1654 ( .o(net_9504), .ck(clk), .d(n8433) );
ms00f80  l1655 ( .o(_net_266), .ck(clk), .d(n8438) );
ms00f80  l1656 ( .o(net_9342), .ck(clk), .d(n8443) );
ms00f80  l1657 ( .o(net_9366), .ck(clk), .d(n8447) );
ms00f80  l1658 ( .o(_net_10477), .ck(clk), .d(n8452) );
ms00f80  l1659 ( .o(net_10388), .ck(clk), .d(n8457) );
ms00f80  l1660 ( .o(net_9587), .ck(clk), .d(n8462) );
ms00f80  l1661 ( .o(_net_128), .ck(clk), .d(n8467) );
ms00f80  l1662 ( .o(_net_9118), .ck(clk), .d(n8472) );
ms00f80  l1663 ( .o(_net_10162), .ck(clk), .d(n8477) );
ms00f80  l1664 ( .o(_net_9382), .ck(clk), .d(n8482) );
ms00f80  l1665 ( .o(net_9486), .ck(clk), .d(n8486) );
ms00f80  l1666 ( .o(_net_231), .ck(clk), .d(n8491) );
ms00f80  l1667 ( .o(net_10006), .ck(clk), .d(n8496) );
ms00f80  l1668 ( .o(net_9443), .ck(clk), .d(n8501) );
ms00f80  l1669 ( .o(net_9433), .ck(clk), .d(n8505) );
ms00f80  l1670 ( .o(_net_9565), .ck(clk), .d(n8510) );
ms00f80  l1671 ( .o(net_108), .ck(clk), .d(n8515) );
ms00f80  l1672 ( .o(net_9655), .ck(clk), .d(n8519) );
ms00f80  l1673 ( .o(_net_10211), .ck(clk), .d(n8524) );
ms00f80  l1674 ( .o(net_9379), .ck(clk), .d(n8529) );
ms00f80  l1675 ( .o(net_9134), .ck(clk), .d(n8534) );
ms00f80  l1676 ( .o(net_9800), .ck(clk), .d(n8538) );
ms00f80  l1677 ( .o(_net_10027), .ck(clk), .d(n8543) );
ms00f80  l1678 ( .o(net_9945), .ck(clk), .d(n8548) );
ms00f80  l1679 ( .o(_net_168), .ck(clk), .d(n8553) );
ms00f80  l1680 ( .o(_net_169), .ck(clk), .d(n8558) );
ms00f80  l1681 ( .o(net_9545), .ck(clk), .d(n8562) );
ms00f80  l1682 ( .o(net_9605), .ck(clk), .d(n8567) );
ms00f80  l1683 ( .o(net_9221), .ck(clk), .d(n8572) );
ms00f80  l1684 ( .o(_net_9117), .ck(clk), .d(n8577) );
ms00f80  l1685 ( .o(net_9621), .ck(clk), .d(n8582) );
ms00f80  l1686 ( .o(net_10064), .ck(clk), .d(n8587) );
ms00f80  l1687 ( .o(_net_9830), .ck(clk), .d(n8592) );
ms00f80  l1688 ( .o(_net_10232), .ck(clk), .d(n8597) );
ms00f80  l1689 ( .o(net_9620), .ck(clk), .d(n8602) );
ms00f80  l1690 ( .o(net_9992), .ck(clk), .d(n8607) );
ms00f80  l1691 ( .o(net_136), .ck(clk), .d(n8612) );
ms00f80  l1692 ( .o(net_225), .ck(clk), .d(n8616) );
ms00f80  l1693 ( .o(_net_9629), .ck(clk), .d(n8621) );
ms00f80  l1694 ( .o(_net_273), .ck(clk), .d(n8626) );
ms00f80  l1695 ( .o(_net_10432), .ck(clk), .d(n8631) );
ms00f80  l1696 ( .o(net_263), .ck(clk), .d(n8636) );
ms00f80  l1697 ( .o(_net_9517), .ck(clk), .d(n8641) );
ms00f80  l1698 ( .o(net_312), .ck(clk), .d(n8646) );
ms00f80  l1699 ( .o(_net_10222), .ck(clk), .d(n8650) );
ms00f80  l1700 ( .o(x1066), .ck(clk), .d(n8655) );
ms00f80  l1701 ( .o(net_9983), .ck(clk), .d(n8659) );
ms00f80  l1702 ( .o(net_9140), .ck(clk), .d(n8664) );
ms00f80  l1703 ( .o(_net_9514), .ck(clk), .d(n8668) );
ms00f80  l1704 ( .o(_net_10406), .ck(clk), .d(n8673) );
ms00f80  l1705 ( .o(net_9995), .ck(clk), .d(n8678) );
ms00f80  l1706 ( .o(net_9825), .ck(clk), .d(n8683) );
ms00f80  l1707 ( .o(_net_9244), .ck(clk), .d(n8688) );
ms00f80  l1708 ( .o(net_9332), .ck(clk), .d(n8693) );
ms00f80  l1709 ( .o(_net_10353), .ck(clk), .d(n8697) );
ms00f80  l1710 ( .o(_net_9315), .ck(clk), .d(n8702) );
ms00f80  l1711 ( .o(_net_10266), .ck(clk), .d(n8707) );
ms00f80  l1712 ( .o(net_192), .ck(clk), .d(n8712) );
ms00f80  l1713 ( .o(_net_10108), .ck(clk), .d(n8717) );
ms00f80  l1714 ( .o(net_10343), .ck(clk), .d(n8722) );
ms00f80  l1715 ( .o(net_9823), .ck(clk), .d(n8727) );
ms00f80  l1716 ( .o(_net_10308), .ck(clk), .d(n8732) );
ms00f80  l1717 ( .o(_net_314), .ck(clk), .d(n8737) );
ms00f80  l1718 ( .o(_net_10154), .ck(clk), .d(n8742) );
ms00f80  l1719 ( .o(_net_10376), .ck(clk), .d(n8747) );
ms00f80  l1720 ( .o(_net_9502), .ck(clk), .d(n8752) );
ms00f80  l1721 ( .o(net_9824), .ck(clk), .d(n8757) );
ms00f80  l1722 ( .o(_net_9630), .ck(clk), .d(n8762) );
ms00f80  l1723 ( .o(_net_10122), .ck(clk), .d(n8767) );
ms00f80  l1724 ( .o(_net_9644), .ck(clk), .d(n8772) );
ms00f80  l1725 ( .o(net_9595), .ck(clk), .d(n8777) );
ms00f80  l1726 ( .o(net_9967), .ck(clk), .d(n8782) );
ms00f80  l1727 ( .o(_net_10365), .ck(clk), .d(n8787) );
ms00f80  l1728 ( .o(net_9146), .ck(clk), .d(n8792) );
ms00f80  l1729 ( .o(net_9871), .ck(clk), .d(n8796) );
ms00f80  l1730 ( .o(x732), .ck(clk), .d(n8800) );
ms00f80  l1731 ( .o(_net_10534), .ck(clk), .d(n8804) );
ms00f80  l1732 ( .o(_net_10167), .ck(clk), .d(n8809) );
ms00f80  l1733 ( .o(net_9662), .ck(clk), .d(n8814) );
ms00f80  l1734 ( .o(net_9717), .ck(clk), .d(n8819) );
ms00f80  l1735 ( .o(net_9955), .ck(clk), .d(n8824) );
ms00f80  l1736 ( .o(_net_9931), .ck(clk), .d(n8829) );
ms00f80  l1737 ( .o(_net_10028), .ck(clk), .d(n8834) );
ms00f80  l1738 ( .o(_net_9735), .ck(clk), .d(n8839) );
ms00f80  l1739 ( .o(_net_10150), .ck(clk), .d(n8844) );
ms00f80  l1740 ( .o(net_9460), .ck(clk), .d(n8849) );
ms00f80  l1741 ( .o(net_9341), .ck(clk), .d(n8853) );
ms00f80  l1742 ( .o(_net_10317), .ck(clk), .d(n8857) );
ms00f80  l1743 ( .o(_net_10223), .ck(clk), .d(n8862) );
ms00f80  l1744 ( .o(_net_10356), .ck(clk), .d(n8867) );
ms00f80  l1745 ( .o(_net_8842), .ck(clk), .d(n8872) );
ms00f80  l1746 ( .o(x1134), .ck(clk), .d(n8876) );

endmodule
